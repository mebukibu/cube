`include "num_data.v"

module w_rom_23 #(
    parameter filename = "../data/data18/weight18_0.txt",
    parameter integer dwidth = `data_len,
    parameter integer awidth = 11,          // 2^11 = 2048 > 5*288 = 1440
    parameter integer words = 5*288
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 18'b000000000100010111;
    mem[1] = 18'b000000000000001001;
    mem[2] = 18'b000000000001101000;
    mem[3] = 18'b111111111111110100;
    mem[4] = 18'b000000000110010110;
    mem[5] = 18'b000000000001111011;
    mem[6] = 18'b000000000110010100;
    mem[7] = 18'b000000000000001011;
    mem[8] = 18'b000000000100100001;
    mem[9] = 18'b111111111011110011;
    mem[10] = 18'b111111001110010011;
    mem[11] = 18'b111111011110101101;
    mem[12] = 18'b111111110101111001;
    mem[13] = 18'b000000000001110111;
    mem[14] = 18'b111111111100010110;
    mem[15] = 18'b000000000001010110;
    mem[16] = 18'b111111011100110001;
    mem[17] = 18'b111111011001110010;
    mem[18] = 18'b111111111101010101;
    mem[19] = 18'b000000000001101001;
    mem[20] = 18'b111111111000001100;
    mem[21] = 18'b000000000000010101;
    mem[22] = 18'b000000000010000100;
    mem[23] = 18'b111111111111000101;
    mem[24] = 18'b000000000001011001;
    mem[25] = 18'b111111111100111110;
    mem[26] = 18'b000000000010101011;
    mem[27] = 18'b111111101010100110;
    mem[28] = 18'b111111011111000101;
    mem[29] = 18'b111111101001001001;
    mem[30] = 18'b111111110100000110;
    mem[31] = 18'b111111100011111101;
    mem[32] = 18'b111111110100011101;
    mem[33] = 18'b000000000001000110;
    mem[34] = 18'b111111111100010100;
    mem[35] = 18'b111111111000011000;
    mem[36] = 18'b000000000000000000;
    mem[37] = 18'b000000000000000000;
    mem[38] = 18'b000000000000000000;
    mem[39] = 18'b000000000000000000;
    mem[40] = 18'b000000000000000000;
    mem[41] = 18'b000000000000000000;
    mem[42] = 18'b000000000000000000;
    mem[43] = 18'b000000000000000000;
    mem[44] = 18'b000000000000000000;
    mem[45] = 18'b000000000000000000;
    mem[46] = 18'b000000000000000000;
    mem[47] = 18'b000000000000000000;
    mem[48] = 18'b000000000000000000;
    mem[49] = 18'b000000000000000000;
    mem[50] = 18'b000000000000000000;
    mem[51] = 18'b000000000000000000;
    mem[52] = 18'b000000000000000000;
    mem[53] = 18'b000000000000000000;
    mem[54] = 18'b000000000000000000;
    mem[55] = 18'b000000000000000000;
    mem[56] = 18'b000000000000000000;
    mem[57] = 18'b000000000000000000;
    mem[58] = 18'b000000000000000000;
    mem[59] = 18'b000000000000000000;
    mem[60] = 18'b000000000000000000;
    mem[61] = 18'b000000000000000000;
    mem[62] = 18'b000000000000000000;
    mem[63] = 18'b000000000000000000;
    mem[64] = 18'b000000000000000000;
    mem[65] = 18'b000000000000000000;
    mem[66] = 18'b000000000000000000;
    mem[67] = 18'b000000000000000000;
    mem[68] = 18'b000000000000000000;
    mem[69] = 18'b000000000000000000;
    mem[70] = 18'b000000000000000000;
    mem[71] = 18'b000000000000000000;
    mem[72] = 18'b000000000000000000;
    mem[73] = 18'b000000000000000000;
    mem[74] = 18'b000000000000000000;
    mem[75] = 18'b000000000000000000;
    mem[76] = 18'b000000000000000000;
    mem[77] = 18'b000000000000000000;
    mem[78] = 18'b000000000000000000;
    mem[79] = 18'b000000000000000000;
    mem[80] = 18'b000000000000000000;
    mem[81] = 18'b000000000000000000;
    mem[82] = 18'b000000000000000000;
    mem[83] = 18'b000000000000000000;
    mem[84] = 18'b000000000000000000;
    mem[85] = 18'b000000000000000000;
    mem[86] = 18'b000000000000000000;
    mem[87] = 18'b000000000000000000;
    mem[88] = 18'b000000000000000000;
    mem[89] = 18'b000000000000000000;
    mem[90] = 18'b000000000000000000;
    mem[91] = 18'b000000000000000000;
    mem[92] = 18'b000000000000000000;
    mem[93] = 18'b000000000000000000;
    mem[94] = 18'b000000000000000000;
    mem[95] = 18'b000000000000000000;
    mem[96] = 18'b000000000000000000;
    mem[97] = 18'b000000000000000000;
    mem[98] = 18'b000000000000000000;
    mem[99] = 18'b000000000000000000;
    mem[100] = 18'b000000000000000000;
    mem[101] = 18'b000000000000000000;
    mem[102] = 18'b000000000000000000;
    mem[103] = 18'b000000000000000000;
    mem[104] = 18'b000000000000000000;
    mem[105] = 18'b000000000000000000;
    mem[106] = 18'b000000000000000000;
    mem[107] = 18'b000000000000000000;
    mem[108] = 18'b000000000000000000;
    mem[109] = 18'b000000000000000000;
    mem[110] = 18'b000000000000000000;
    mem[111] = 18'b000000000000000000;
    mem[112] = 18'b000000000000000000;
    mem[113] = 18'b000000000000000000;
    mem[114] = 18'b000000000000000000;
    mem[115] = 18'b000000000000000000;
    mem[116] = 18'b000000000000000000;
    mem[117] = 18'b000000000000000000;
    mem[118] = 18'b000000000000000000;
    mem[119] = 18'b000000000000000000;
    mem[120] = 18'b000000000000000000;
    mem[121] = 18'b000000000000000000;
    mem[122] = 18'b000000000000000000;
    mem[123] = 18'b000000000000000000;
    mem[124] = 18'b000000000000000000;
    mem[125] = 18'b000000000000000000;
    mem[126] = 18'b000000000000000000;
    mem[127] = 18'b000000000000000000;
    mem[128] = 18'b000000000000000000;
    mem[129] = 18'b000000000000000000;
    mem[130] = 18'b000000000000000000;
    mem[131] = 18'b000000000000000000;
    mem[132] = 18'b000000000000000000;
    mem[133] = 18'b000000000000000000;
    mem[134] = 18'b000000000000000000;
    mem[135] = 18'b000000000000000000;
    mem[136] = 18'b000000000000000000;
    mem[137] = 18'b000000000000000000;
    mem[138] = 18'b000000000000000000;
    mem[139] = 18'b000000000000000000;
    mem[140] = 18'b000000000000000000;
    mem[141] = 18'b000000000000000000;
    mem[142] = 18'b000000000000000000;
    mem[143] = 18'b000000000000000000;
    mem[144] = 18'b000000000000000000;
    mem[145] = 18'b000000000000000000;
    mem[146] = 18'b000000000000000000;
    mem[147] = 18'b000000000000000000;
    mem[148] = 18'b000000000000000000;
    mem[149] = 18'b000000000000000000;
    mem[150] = 18'b000000000000000000;
    mem[151] = 18'b000000000000000000;
    mem[152] = 18'b000000000000000000;
    mem[153] = 18'b000000000000000000;
    mem[154] = 18'b000000000000000000;
    mem[155] = 18'b000000000000000000;
    mem[156] = 18'b000000000000000000;
    mem[157] = 18'b000000000000000000;
    mem[158] = 18'b000000000000000000;
    mem[159] = 18'b000000000000000000;
    mem[160] = 18'b000000000000000000;
    mem[161] = 18'b000000000000000000;
    mem[162] = 18'b000000000000000000;
    mem[163] = 18'b000000000000000000;
    mem[164] = 18'b000000000000000000;
    mem[165] = 18'b000000000000000000;
    mem[166] = 18'b000000000000000000;
    mem[167] = 18'b000000000000000000;
    mem[168] = 18'b000000000000000000;
    mem[169] = 18'b000000000000000000;
    mem[170] = 18'b000000000000000000;
    mem[171] = 18'b000000000000000000;
    mem[172] = 18'b000000000000000000;
    mem[173] = 18'b000000000000000000;
    mem[174] = 18'b000000000000000000;
    mem[175] = 18'b000000000000000000;
    mem[176] = 18'b000000000000000000;
    mem[177] = 18'b000000000000000000;
    mem[178] = 18'b000000000000000000;
    mem[179] = 18'b000000000000000000;
    mem[180] = 18'b000000000000000000;
    mem[181] = 18'b000000000000000000;
    mem[182] = 18'b000000000000000000;
    mem[183] = 18'b000000000000000000;
    mem[184] = 18'b000000000000000000;
    mem[185] = 18'b000000000000000000;
    mem[186] = 18'b000000000000000000;
    mem[187] = 18'b000000000000000000;
    mem[188] = 18'b000000000000000000;
    mem[189] = 18'b000000000000000000;
    mem[190] = 18'b000000000000000000;
    mem[191] = 18'b000000000000000000;
    mem[192] = 18'b000000000000000000;
    mem[193] = 18'b000000000000000000;
    mem[194] = 18'b000000000000000000;
    mem[195] = 18'b000000000000000000;
    mem[196] = 18'b000000000000000000;
    mem[197] = 18'b000000000000000000;
    mem[198] = 18'b000000000000000000;
    mem[199] = 18'b000000000000000000;
    mem[200] = 18'b000000000000000000;
    mem[201] = 18'b000000000000000000;
    mem[202] = 18'b000000000000000000;
    mem[203] = 18'b000000000000000000;
    mem[204] = 18'b000000000000000000;
    mem[205] = 18'b000000000000000000;
    mem[206] = 18'b000000000000000000;
    mem[207] = 18'b000000000000000000;
    mem[208] = 18'b000000000000000000;
    mem[209] = 18'b000000000000000000;
    mem[210] = 18'b000000000000000000;
    mem[211] = 18'b000000000000000000;
    mem[212] = 18'b000000000000000000;
    mem[213] = 18'b000000000000000000;
    mem[214] = 18'b000000000000000000;
    mem[215] = 18'b000000000000000000;
    mem[216] = 18'b000000000000000000;
    mem[217] = 18'b000000000000000000;
    mem[218] = 18'b000000000000000000;
    mem[219] = 18'b000000000000000000;
    mem[220] = 18'b000000000000000000;
    mem[221] = 18'b000000000000000000;
    mem[222] = 18'b000000000000000000;
    mem[223] = 18'b000000000000000000;
    mem[224] = 18'b000000000000000000;
    mem[225] = 18'b000000000000000000;
    mem[226] = 18'b000000000000000000;
    mem[227] = 18'b000000000000000000;
    mem[228] = 18'b000000000000000000;
    mem[229] = 18'b000000000000000000;
    mem[230] = 18'b000000000000000000;
    mem[231] = 18'b000000000000000000;
    mem[232] = 18'b000000000000000000;
    mem[233] = 18'b000000000000000000;
    mem[234] = 18'b000000000000000000;
    mem[235] = 18'b000000000000000000;
    mem[236] = 18'b000000000000000000;
    mem[237] = 18'b000000000000000000;
    mem[238] = 18'b000000000000000000;
    mem[239] = 18'b000000000000000000;
    mem[240] = 18'b000000000000000000;
    mem[241] = 18'b000000000000000000;
    mem[242] = 18'b000000000000000000;
    mem[243] = 18'b000000000000000000;
    mem[244] = 18'b000000000000000000;
    mem[245] = 18'b000000000000000000;
    mem[246] = 18'b000000000000000000;
    mem[247] = 18'b000000000000000000;
    mem[248] = 18'b000000000000000000;
    mem[249] = 18'b000000000000000000;
    mem[250] = 18'b000000000000000000;
    mem[251] = 18'b000000000000000000;
    mem[252] = 18'b000000000000000000;
    mem[253] = 18'b000000000000000000;
    mem[254] = 18'b000000000000000000;
    mem[255] = 18'b000000000000000000;
    mem[256] = 18'b000000000000000000;
    mem[257] = 18'b000000000000000000;
    mem[258] = 18'b000000000000000000;
    mem[259] = 18'b000000000000000000;
    mem[260] = 18'b000000000000000000;
    mem[261] = 18'b000000000000000000;
    mem[262] = 18'b000000000000000000;
    mem[263] = 18'b000000000000000000;
    mem[264] = 18'b000000000000000000;
    mem[265] = 18'b000000000000000000;
    mem[266] = 18'b000000000000000000;
    mem[267] = 18'b000000000000000000;
    mem[268] = 18'b000000000000000000;
    mem[269] = 18'b000000000000000000;
    mem[270] = 18'b000000000000000000;
    mem[271] = 18'b000000000000000000;
    mem[272] = 18'b000000000000000000;
    mem[273] = 18'b000000000000000000;
    mem[274] = 18'b000000000000000000;
    mem[275] = 18'b000000000000000000;
    mem[276] = 18'b000000000000000000;
    mem[277] = 18'b000000000000000000;
    mem[278] = 18'b000000000000000000;
    mem[279] = 18'b000000000000000000;
    mem[280] = 18'b000000000000000000;
    mem[281] = 18'b000000000000000000;
    mem[282] = 18'b000000000000000000;
    mem[283] = 18'b000000000000000000;
    mem[284] = 18'b000000000000000000;
    mem[285] = 18'b000000000000000000;
    mem[286] = 18'b000000000000000000;
    mem[287] = 18'b000000000000000000;
    mem[288] = 18'b111111111100111110;
    mem[289] = 18'b111111110110011001;
    mem[290] = 18'b111111110111000010;
    mem[291] = 18'b111111111110111001;
    mem[292] = 18'b000000000011110100;
    mem[293] = 18'b000000000000111100;
    mem[294] = 18'b111111111100000001;
    mem[295] = 18'b000000000110101101;
    mem[296] = 18'b111111110101010001;
    mem[297] = 18'b111111111100000111;
    mem[298] = 18'b111111111000111100;
    mem[299] = 18'b111111111010111010;
    mem[300] = 18'b111111111110110100;
    mem[301] = 18'b000000000101101101;
    mem[302] = 18'b111111111111111101;
    mem[303] = 18'b000000000111010000;
    mem[304] = 18'b000000000100101000;
    mem[305] = 18'b000000000011110101;
    mem[306] = 18'b000000000111000001;
    mem[307] = 18'b111111111100110111;
    mem[308] = 18'b111111111001001111;
    mem[309] = 18'b111111111011001110;
    mem[310] = 18'b111111111101001101;
    mem[311] = 18'b000000000001001100;
    mem[312] = 18'b000000000001001100;
    mem[313] = 18'b000000000110000011;
    mem[314] = 18'b000000000011110001;
    mem[315] = 18'b000000000010010100;
    mem[316] = 18'b111111111100010110;
    mem[317] = 18'b111111111011001110;
    mem[318] = 18'b000000000110111100;
    mem[319] = 18'b111111111110001111;
    mem[320] = 18'b000000000110010011;
    mem[321] = 18'b111111111010000011;
    mem[322] = 18'b111111111111110100;
    mem[323] = 18'b111111111101111001;
    mem[324] = 18'b000000000100110101;
    mem[325] = 18'b111111111101010000;
    mem[326] = 18'b000000000111110101;
    mem[327] = 18'b111111111110100101;
    mem[328] = 18'b000000000000011110;
    mem[329] = 18'b000000000010001011;
    mem[330] = 18'b000000001000001111;
    mem[331] = 18'b111111111101110000;
    mem[332] = 18'b000000000101011101;
    mem[333] = 18'b111111111101001000;
    mem[334] = 18'b111111111110010100;
    mem[335] = 18'b000000000001101011;
    mem[336] = 18'b111111111101001000;
    mem[337] = 18'b111111111110111101;
    mem[338] = 18'b000000000100011011;
    mem[339] = 18'b000000000010111011;
    mem[340] = 18'b000000000010101000;
    mem[341] = 18'b111111111101101101;
    mem[342] = 18'b111111111101100110;
    mem[343] = 18'b000000000100001001;
    mem[344] = 18'b000000000100101101;
    mem[345] = 18'b000000001010110111;
    mem[346] = 18'b000000000001110110;
    mem[347] = 18'b000000000010110000;
    mem[348] = 18'b000000000011011110;
    mem[349] = 18'b000000000001111011;
    mem[350] = 18'b000000001000000010;
    mem[351] = 18'b111111111101000111;
    mem[352] = 18'b111111111011100000;
    mem[353] = 18'b111111111110101110;
    mem[354] = 18'b000000000100000001;
    mem[355] = 18'b000000000000001101;
    mem[356] = 18'b111111111110011001;
    mem[357] = 18'b111111111100101011;
    mem[358] = 18'b000000000100010111;
    mem[359] = 18'b111111111111001000;
    mem[360] = 18'b000000000011110101;
    mem[361] = 18'b111111111011000101;
    mem[362] = 18'b000000000011111100;
    mem[363] = 18'b000000000001010101;
    mem[364] = 18'b111111111101100001;
    mem[365] = 18'b000000000010010110;
    mem[366] = 18'b000000000010011111;
    mem[367] = 18'b000000000111000100;
    mem[368] = 18'b000000000000111100;
    mem[369] = 18'b111111111010101000;
    mem[370] = 18'b111111111100100000;
    mem[371] = 18'b000000000000110011;
    mem[372] = 18'b000000001001101101;
    mem[373] = 18'b111111110101011111;
    mem[374] = 18'b000000000110011000;
    mem[375] = 18'b000000000011100100;
    mem[376] = 18'b111111111000110000;
    mem[377] = 18'b111111111011000000;
    mem[378] = 18'b000000000010111100;
    mem[379] = 18'b000000000000110000;
    mem[380] = 18'b111111111101001011;
    mem[381] = 18'b000000000101011000;
    mem[382] = 18'b111111111100010010;
    mem[383] = 18'b111111111100010010;
    mem[384] = 18'b000000001010000100;
    mem[385] = 18'b000000000000111100;
    mem[386] = 18'b000000001001001010;
    mem[387] = 18'b111111111010000011;
    mem[388] = 18'b000000000010001111;
    mem[389] = 18'b000000000011011011;
    mem[390] = 18'b000000000100000100;
    mem[391] = 18'b000000000001011111;
    mem[392] = 18'b000000010000100110;
    mem[393] = 18'b111111111101100010;
    mem[394] = 18'b000000000011010010;
    mem[395] = 18'b000000001001001110;
    mem[396] = 18'b111111111110000011;
    mem[397] = 18'b111111111100101010;
    mem[398] = 18'b000000000100010010;
    mem[399] = 18'b111111111111101000;
    mem[400] = 18'b000000000001111000;
    mem[401] = 18'b111111111111001100;
    mem[402] = 18'b111111111001010110;
    mem[403] = 18'b000000000100000111;
    mem[404] = 18'b111111111100111010;
    mem[405] = 18'b111111111001101010;
    mem[406] = 18'b000000000010011011;
    mem[407] = 18'b111111111010011110;
    mem[408] = 18'b111111111011111001;
    mem[409] = 18'b000000000000101100;
    mem[410] = 18'b111111110100100101;
    mem[411] = 18'b111111111011101111;
    mem[412] = 18'b000000000001001110;
    mem[413] = 18'b111111111111101010;
    mem[414] = 18'b111111110110110010;
    mem[415] = 18'b111111111011101010;
    mem[416] = 18'b000000000100010001;
    mem[417] = 18'b111111111110011001;
    mem[418] = 18'b111111111111110011;
    mem[419] = 18'b111111110110001111;
    mem[420] = 18'b111111110111111111;
    mem[421] = 18'b000000000010110000;
    mem[422] = 18'b000000001010100000;
    mem[423] = 18'b111111111111100010;
    mem[424] = 18'b000000000100010000;
    mem[425] = 18'b000000000100011100;
    mem[426] = 18'b111111111111110001;
    mem[427] = 18'b111111111011111110;
    mem[428] = 18'b111111110111010001;
    mem[429] = 18'b111111111101110101;
    mem[430] = 18'b000000000000011111;
    mem[431] = 18'b000000000111100100;
    mem[432] = 18'b000000000001100001;
    mem[433] = 18'b111111111111110110;
    mem[434] = 18'b111111110101110001;
    mem[435] = 18'b000000000101011101;
    mem[436] = 18'b000000000011011100;
    mem[437] = 18'b111111111110010011;
    mem[438] = 18'b111111111110010111;
    mem[439] = 18'b111111110011010000;
    mem[440] = 18'b111111111110010000;
    mem[441] = 18'b111111111100000011;
    mem[442] = 18'b000000000010101100;
    mem[443] = 18'b000000001000001111;
    mem[444] = 18'b111111111000011000;
    mem[445] = 18'b111111111001011101;
    mem[446] = 18'b000000000001111001;
    mem[447] = 18'b111111111011000101;
    mem[448] = 18'b111111111111000110;
    mem[449] = 18'b000000000101001011;
    mem[450] = 18'b111111111001110111;
    mem[451] = 18'b111111111011111011;
    mem[452] = 18'b000000000101100011;
    mem[453] = 18'b111111111110111001;
    mem[454] = 18'b111111111111100101;
    mem[455] = 18'b111111111001101011;
    mem[456] = 18'b111111111011000101;
    mem[457] = 18'b000000000111000011;
    mem[458] = 18'b000000001010111000;
    mem[459] = 18'b000000000111010011;
    mem[460] = 18'b000000000001001010;
    mem[461] = 18'b111111111110100010;
    mem[462] = 18'b000000000111011011;
    mem[463] = 18'b111111111111101001;
    mem[464] = 18'b000000000011001100;
    mem[465] = 18'b000000000110001010;
    mem[466] = 18'b000000000101100001;
    mem[467] = 18'b000000000010100111;
    mem[468] = 18'b000000000001100011;
    mem[469] = 18'b111111111100010101;
    mem[470] = 18'b111111111011001111;
    mem[471] = 18'b000000000001101101;
    mem[472] = 18'b000000000010011110;
    mem[473] = 18'b000000000110010110;
    mem[474] = 18'b000000000110111001;
    mem[475] = 18'b000000000101001000;
    mem[476] = 18'b000000000001101001;
    mem[477] = 18'b000000000000010001;
    mem[478] = 18'b111111111011010110;
    mem[479] = 18'b111111111110001101;
    mem[480] = 18'b000000000100000100;
    mem[481] = 18'b111111111101111011;
    mem[482] = 18'b111111111110010010;
    mem[483] = 18'b111111111001100111;
    mem[484] = 18'b000000001000111010;
    mem[485] = 18'b000000000100110011;
    mem[486] = 18'b000000000001000111;
    mem[487] = 18'b111111111110001001;
    mem[488] = 18'b000000000011100011;
    mem[489] = 18'b111111111111111010;
    mem[490] = 18'b000000000101111101;
    mem[491] = 18'b111111111101000101;
    mem[492] = 18'b111111111001011001;
    mem[493] = 18'b111111111101110011;
    mem[494] = 18'b111111111110010011;
    mem[495] = 18'b000000000111100100;
    mem[496] = 18'b111111111101110111;
    mem[497] = 18'b111111111100001111;
    mem[498] = 18'b000000000001111111;
    mem[499] = 18'b111111111101101100;
    mem[500] = 18'b111111111111001010;
    mem[501] = 18'b111111111101011111;
    mem[502] = 18'b000000000100001011;
    mem[503] = 18'b000000000011011001;
    mem[504] = 18'b111111111111001001;
    mem[505] = 18'b000000000011011011;
    mem[506] = 18'b111111111010011001;
    mem[507] = 18'b000000001000111011;
    mem[508] = 18'b111111110111101000;
    mem[509] = 18'b111111111111001000;
    mem[510] = 18'b111111110111011010;
    mem[511] = 18'b000000000011010110;
    mem[512] = 18'b111111111100100110;
    mem[513] = 18'b111111111111001011;
    mem[514] = 18'b111111111111010111;
    mem[515] = 18'b111111111010110011;
    mem[516] = 18'b111111111111010100;
    mem[517] = 18'b000000000011111000;
    mem[518] = 18'b000000000010100001;
    mem[519] = 18'b000000000010111110;
    mem[520] = 18'b000000000011101010;
    mem[521] = 18'b000000000001010001;
    mem[522] = 18'b000000000010101110;
    mem[523] = 18'b000000000000001111;
    mem[524] = 18'b111111111100010001;
    mem[525] = 18'b000000000101101100;
    mem[526] = 18'b000000000101111011;
    mem[527] = 18'b111111111110111001;
    mem[528] = 18'b000000000110000100;
    mem[529] = 18'b111111111110111010;
    mem[530] = 18'b000000000100010000;
    mem[531] = 18'b000000000000001000;
    mem[532] = 18'b000000000101001010;
    mem[533] = 18'b111111111111101011;
    mem[534] = 18'b000000000111100110;
    mem[535] = 18'b111111111101100011;
    mem[536] = 18'b111111111101100011;
    mem[537] = 18'b111111111001110110;
    mem[538] = 18'b000000000001110101;
    mem[539] = 18'b000000000010001110;
    mem[540] = 18'b111111111101101000;
    mem[541] = 18'b000000001000000011;
    mem[542] = 18'b000000000001110111;
    mem[543] = 18'b111111111000111110;
    mem[544] = 18'b111111111111001111;
    mem[545] = 18'b000000000110110010;
    mem[546] = 18'b000000000000100111;
    mem[547] = 18'b000000000000010101;
    mem[548] = 18'b000000000001110011;
    mem[549] = 18'b111111110101101011;
    mem[550] = 18'b111111111101000011;
    mem[551] = 18'b111111111110011011;
    mem[552] = 18'b111111111110111011;
    mem[553] = 18'b111111111101001010;
    mem[554] = 18'b111111111100011111;
    mem[555] = 18'b000000000111010010;
    mem[556] = 18'b000000000101001110;
    mem[557] = 18'b000000000001110000;
    mem[558] = 18'b111111111100100111;
    mem[559] = 18'b000000000001101000;
    mem[560] = 18'b000000000110010110;
    mem[561] = 18'b111111111110110001;
    mem[562] = 18'b111111111111010010;
    mem[563] = 18'b000000000111010001;
    mem[564] = 18'b111111111010110110;
    mem[565] = 18'b111111111011101000;
    mem[566] = 18'b111111111011100100;
    mem[567] = 18'b000000000100110010;
    mem[568] = 18'b000000000010011110;
    mem[569] = 18'b000000000101101100;
    mem[570] = 18'b000000000010110101;
    mem[571] = 18'b000000000010000100;
    mem[572] = 18'b000000000001100000;
    mem[573] = 18'b111111111101010001;
    mem[574] = 18'b111111111100101101;
    mem[575] = 18'b000000000001000111;
    mem[576] = 18'b000000000000011100;
    mem[577] = 18'b000000000010000100;
    mem[578] = 18'b111111111110011010;
    mem[579] = 18'b111111111110101000;
    mem[580] = 18'b000000000011100101;
    mem[581] = 18'b111111111100101111;
    mem[582] = 18'b000000000100000001;
    mem[583] = 18'b000000000010000010;
    mem[584] = 18'b111111111111000010;
    mem[585] = 18'b000000000001100101;
    mem[586] = 18'b000000000101000111;
    mem[587] = 18'b000000000100000101;
    mem[588] = 18'b000000000000100100;
    mem[589] = 18'b111111111011000011;
    mem[590] = 18'b111111111001111101;
    mem[591] = 18'b111111111000111111;
    mem[592] = 18'b111111111111111010;
    mem[593] = 18'b111111111101111110;
    mem[594] = 18'b000000000001101011;
    mem[595] = 18'b111111111100100110;
    mem[596] = 18'b000000000101001100;
    mem[597] = 18'b111111111111010110;
    mem[598] = 18'b111111111011100110;
    mem[599] = 18'b000000000000100111;
    mem[600] = 18'b111111111100101100;
    mem[601] = 18'b000000000010101111;
    mem[602] = 18'b000000000001010000;
    mem[603] = 18'b000000000010111001;
    mem[604] = 18'b000000000001101101;
    mem[605] = 18'b111111111110100110;
    mem[606] = 18'b000000000000010001;
    mem[607] = 18'b111111111100111100;
    mem[608] = 18'b111111111001000011;
    mem[609] = 18'b000000000100110001;
    mem[610] = 18'b111111111111000011;
    mem[611] = 18'b000000000100000010;
    mem[612] = 18'b111111111101001110;
    mem[613] = 18'b000000000000000111;
    mem[614] = 18'b111111111010111000;
    mem[615] = 18'b111111111100110101;
    mem[616] = 18'b000000000010001100;
    mem[617] = 18'b111111111010000000;
    mem[618] = 18'b000000000111001001;
    mem[619] = 18'b000000000000000000;
    mem[620] = 18'b111111110111001111;
    mem[621] = 18'b000000000000100000;
    mem[622] = 18'b000000000111000010;
    mem[623] = 18'b000000000011010110;
    mem[624] = 18'b000000000001010011;
    mem[625] = 18'b000000000000001011;
    mem[626] = 18'b111111111001101100;
    mem[627] = 18'b111111111111111011;
    mem[628] = 18'b111111111111000111;
    mem[629] = 18'b111111111001101101;
    mem[630] = 18'b111111111011101010;
    mem[631] = 18'b000000000001111110;
    mem[632] = 18'b000000000001001001;
    mem[633] = 18'b111111111110000100;
    mem[634] = 18'b000000000000101100;
    mem[635] = 18'b000000000110101011;
    mem[636] = 18'b000000000111011000;
    mem[637] = 18'b111111111100110001;
    mem[638] = 18'b000000000000111011;
    mem[639] = 18'b111111111100101010;
    mem[640] = 18'b111111111011001100;
    mem[641] = 18'b000000000011010001;
    mem[642] = 18'b111111111111101000;
    mem[643] = 18'b111111111111111011;
    mem[644] = 18'b111111111111100000;
    mem[645] = 18'b000000000000111111;
    mem[646] = 18'b111111111101100001;
    mem[647] = 18'b000000000000011000;
    mem[648] = 18'b111111111111011001;
    mem[649] = 18'b111111111111100100;
    mem[650] = 18'b111111111101101111;
    mem[651] = 18'b111111111011111001;
    mem[652] = 18'b111111111010011011;
    mem[653] = 18'b111111111111011101;
    mem[654] = 18'b000000000011101001;
    mem[655] = 18'b111111111110000011;
    mem[656] = 18'b111111111111110110;
    mem[657] = 18'b111111111100001001;
    mem[658] = 18'b000000000010001010;
    mem[659] = 18'b000000000101101010;
    mem[660] = 18'b111111111111010100;
    mem[661] = 18'b111111111110011000;
    mem[662] = 18'b000000000010010110;
    mem[663] = 18'b000000000000101000;
    mem[664] = 18'b111111111101000111;
    mem[665] = 18'b000000000000110100;
    mem[666] = 18'b111111111101110101;
    mem[667] = 18'b000000001000000011;
    mem[668] = 18'b111111111100101110;
    mem[669] = 18'b111111111001011000;
    mem[670] = 18'b111111111110010001;
    mem[671] = 18'b000000000010000001;
    mem[672] = 18'b111111111110100101;
    mem[673] = 18'b000000000000110010;
    mem[674] = 18'b111111111101011011;
    mem[675] = 18'b111111111000011111;
    mem[676] = 18'b000000000011010110;
    mem[677] = 18'b111111111101110111;
    mem[678] = 18'b111111111111100110;
    mem[679] = 18'b000000000010010011;
    mem[680] = 18'b000000000000111101;
    mem[681] = 18'b000000000100001000;
    mem[682] = 18'b000000000011100111;
    mem[683] = 18'b000000000000110000;
    mem[684] = 18'b000000000110011110;
    mem[685] = 18'b000000000111000001;
    mem[686] = 18'b000000000110100011;
    mem[687] = 18'b111111111111010011;
    mem[688] = 18'b000000000101101001;
    mem[689] = 18'b000000000100000100;
    mem[690] = 18'b000000000010110111;
    mem[691] = 18'b000000000111001101;
    mem[692] = 18'b000000000100010011;
    mem[693] = 18'b111111111111110100;
    mem[694] = 18'b111111111001100011;
    mem[695] = 18'b111111111000000001;
    mem[696] = 18'b000000000001000100;
    mem[697] = 18'b111111111011110111;
    mem[698] = 18'b111111111110110011;
    mem[699] = 18'b111111111101001101;
    mem[700] = 18'b000000001000010100;
    mem[701] = 18'b000000001000110001;
    mem[702] = 18'b000000000001001001;
    mem[703] = 18'b000000000110001100;
    mem[704] = 18'b000000000101100101;
    mem[705] = 18'b111111111011110101;
    mem[706] = 18'b111111111110011001;
    mem[707] = 18'b000000001010001100;
    mem[708] = 18'b000000000101111001;
    mem[709] = 18'b000000000101010001;
    mem[710] = 18'b000000000101110100;
    mem[711] = 18'b000000000010101001;
    mem[712] = 18'b111111111111110110;
    mem[713] = 18'b000000000000001000;
    mem[714] = 18'b111111111110100110;
    mem[715] = 18'b000000000101101100;
    mem[716] = 18'b000000000001100111;
    mem[717] = 18'b111111111010101111;
    mem[718] = 18'b111111111111100000;
    mem[719] = 18'b000000000010000110;
    mem[720] = 18'b000000000011010111;
    mem[721] = 18'b000000000010011100;
    mem[722] = 18'b000000000000011010;
    mem[723] = 18'b111111111001101010;
    mem[724] = 18'b111111111110000000;
    mem[725] = 18'b111111111101011010;
    mem[726] = 18'b000000000110000000;
    mem[727] = 18'b000000000111110110;
    mem[728] = 18'b111111111010001000;
    mem[729] = 18'b111111111111100010;
    mem[730] = 18'b111111111001011101;
    mem[731] = 18'b000000000000101110;
    mem[732] = 18'b111111111110000111;
    mem[733] = 18'b111111111100010001;
    mem[734] = 18'b111111111011110110;
    mem[735] = 18'b111111111111011000;
    mem[736] = 18'b111111110111111101;
    mem[737] = 18'b000000000001100001;
    mem[738] = 18'b000000000011110110;
    mem[739] = 18'b000000000000111110;
    mem[740] = 18'b000000000010001110;
    mem[741] = 18'b000000000101011111;
    mem[742] = 18'b111111111100000101;
    mem[743] = 18'b111111111110110010;
    mem[744] = 18'b000000000001111100;
    mem[745] = 18'b111111111011110001;
    mem[746] = 18'b000000000001011110;
    mem[747] = 18'b111111111111101101;
    mem[748] = 18'b000000000011011001;
    mem[749] = 18'b000000000100001010;
    mem[750] = 18'b111111111101001011;
    mem[751] = 18'b000000001000011110;
    mem[752] = 18'b111111111010111111;
    mem[753] = 18'b000000000000011101;
    mem[754] = 18'b000000000100011110;
    mem[755] = 18'b111111111110010110;
    mem[756] = 18'b111111111111001100;
    mem[757] = 18'b111111111100011001;
    mem[758] = 18'b000000000011001000;
    mem[759] = 18'b111111111101001010;
    mem[760] = 18'b111111111100101101;
    mem[761] = 18'b000000000001001101;
    mem[762] = 18'b111111111011000100;
    mem[763] = 18'b111111111010011000;
    mem[764] = 18'b000000000100110101;
    mem[765] = 18'b111111111111100001;
    mem[766] = 18'b111111111111101110;
    mem[767] = 18'b000000000011111011;
    mem[768] = 18'b000000000011101000;
    mem[769] = 18'b111111111011010011;
    mem[770] = 18'b111111111110101011;
    mem[771] = 18'b111111111100101000;
    mem[772] = 18'b111111111110010100;
    mem[773] = 18'b111111111110111100;
    mem[774] = 18'b000000000111111000;
    mem[775] = 18'b000000001100111011;
    mem[776] = 18'b000000001110100111;
    mem[777] = 18'b000000000001010011;
    mem[778] = 18'b000000000011001111;
    mem[779] = 18'b000000000110011100;
    mem[780] = 18'b000000000110010110;
    mem[781] = 18'b000000000111011011;
    mem[782] = 18'b000000000011011110;
    mem[783] = 18'b111111111111011010;
    mem[784] = 18'b000000000000101110;
    mem[785] = 18'b111111111011010100;
    mem[786] = 18'b000000000001000010;
    mem[787] = 18'b000000000010010100;
    mem[788] = 18'b000000000100100011;
    mem[789] = 18'b111111111101000001;
    mem[790] = 18'b000000000011000000;
    mem[791] = 18'b111111111101101101;
    mem[792] = 18'b111111111010001100;
    mem[793] = 18'b000000000000111100;
    mem[794] = 18'b111111111001011000;
    mem[795] = 18'b111111111110001001;
    mem[796] = 18'b111111111101010000;
    mem[797] = 18'b000000000000010011;
    mem[798] = 18'b111111111110110000;
    mem[799] = 18'b000000000001011000;
    mem[800] = 18'b000000000001000000;
    mem[801] = 18'b111111111110011111;
    mem[802] = 18'b111111111100011110;
    mem[803] = 18'b111111111111110110;
    mem[804] = 18'b000000000100010011;
    mem[805] = 18'b111111111110101000;
    mem[806] = 18'b111111111111100111;
    mem[807] = 18'b111111111101000011;
    mem[808] = 18'b000000000000110010;
    mem[809] = 18'b111111111010111111;
    mem[810] = 18'b111111111011001100;
    mem[811] = 18'b000000000010011111;
    mem[812] = 18'b111111111101110001;
    mem[813] = 18'b000000000001110110;
    mem[814] = 18'b111111111111111100;
    mem[815] = 18'b111111111001110111;
    mem[816] = 18'b000000000101111101;
    mem[817] = 18'b000000000010110001;
    mem[818] = 18'b111111111101011100;
    mem[819] = 18'b000000000001110110;
    mem[820] = 18'b000000001000011110;
    mem[821] = 18'b000000000101010111;
    mem[822] = 18'b000000000010100010;
    mem[823] = 18'b000000000000110001;
    mem[824] = 18'b000000000100011111;
    mem[825] = 18'b000000000101001101;
    mem[826] = 18'b000000000000101011;
    mem[827] = 18'b111111110101100110;
    mem[828] = 18'b111111111111000001;
    mem[829] = 18'b111111111000111100;
    mem[830] = 18'b000000000011100011;
    mem[831] = 18'b111111111100110001;
    mem[832] = 18'b000000000000011100;
    mem[833] = 18'b000000000001010000;
    mem[834] = 18'b111111111110101100;
    mem[835] = 18'b111111111111011000;
    mem[836] = 18'b000000000100111000;
    mem[837] = 18'b000000000101000101;
    mem[838] = 18'b111111111110000010;
    mem[839] = 18'b000000000010100001;
    mem[840] = 18'b111111111110100001;
    mem[841] = 18'b000000000000001100;
    mem[842] = 18'b111111111111011001;
    mem[843] = 18'b111111111100101110;
    mem[844] = 18'b111111111001000011;
    mem[845] = 18'b000000000000100111;
    mem[846] = 18'b111111111101011101;
    mem[847] = 18'b111111111011010000;
    mem[848] = 18'b000000000000100101;
    mem[849] = 18'b111111111011011011;
    mem[850] = 18'b111111111111010011;
    mem[851] = 18'b000000000000011111;
    mem[852] = 18'b000000000010011000;
    mem[853] = 18'b111111111110101011;
    mem[854] = 18'b111111111010011010;
    mem[855] = 18'b000000000000001000;
    mem[856] = 18'b000000000110001111;
    mem[857] = 18'b000000000100110111;
    mem[858] = 18'b111111111111100101;
    mem[859] = 18'b111111111101001101;
    mem[860] = 18'b111111111111001111;
    mem[861] = 18'b111111110110100010;
    mem[862] = 18'b000000000001000011;
    mem[863] = 18'b111111111101101001;
    mem[864] = 18'b111111111111111010;
    mem[865] = 18'b000000000000000001;
    mem[866] = 18'b000000000000000100;
    mem[867] = 18'b000000000000011001;
    mem[868] = 18'b000000000000011110;
    mem[869] = 18'b111111111111100011;
    mem[870] = 18'b111111111111111101;
    mem[871] = 18'b000000000000001111;
    mem[872] = 18'b000000000000000100;
    mem[873] = 18'b000000000000001111;
    mem[874] = 18'b111111111111110111;
    mem[875] = 18'b111111111111100000;
    mem[876] = 18'b111111111111110101;
    mem[877] = 18'b111111111111111101;
    mem[878] = 18'b000000000000010010;
    mem[879] = 18'b000000000000010010;
    mem[880] = 18'b000000000000000101;
    mem[881] = 18'b111111111111110001;
    mem[882] = 18'b000000000000000111;
    mem[883] = 18'b000000000000001000;
    mem[884] = 18'b000000000000000101;
    mem[885] = 18'b111111111111111001;
    mem[886] = 18'b000000000000011101;
    mem[887] = 18'b111111111111111101;
    mem[888] = 18'b000000000000101010;
    mem[889] = 18'b000000000000000100;
    mem[890] = 18'b000000000000010101;
    mem[891] = 18'b111111111111110100;
    mem[892] = 18'b111111111111110011;
    mem[893] = 18'b111111111111110110;
    mem[894] = 18'b000000000000001011;
    mem[895] = 18'b111111111111110111;
    mem[896] = 18'b111111111111101001;
    mem[897] = 18'b000000000000011110;
    mem[898] = 18'b000000000000001101;
    mem[899] = 18'b111111111111111010;
    mem[900] = 18'b000000000000000100;
    mem[901] = 18'b000000000000001010;
    mem[902] = 18'b000000000000001100;
    mem[903] = 18'b000000000000000100;
    mem[904] = 18'b000000000000001111;
    mem[905] = 18'b000000000000010001;
    mem[906] = 18'b000000000000000111;
    mem[907] = 18'b000000000000001011;
    mem[908] = 18'b000000000000100010;
    mem[909] = 18'b000000000000011110;
    mem[910] = 18'b000000000000000011;
    mem[911] = 18'b000000000000001000;
    mem[912] = 18'b111111111111110000;
    mem[913] = 18'b000000000000010000;
    mem[914] = 18'b000000000000001001;
    mem[915] = 18'b000000000000010010;
    mem[916] = 18'b111111111111110001;
    mem[917] = 18'b111111111111100001;
    mem[918] = 18'b111111111111111110;
    mem[919] = 18'b000000000000010001;
    mem[920] = 18'b000000000000010010;
    mem[921] = 18'b000000000000010011;
    mem[922] = 18'b000000000000010000;
    mem[923] = 18'b000000000000010100;
    mem[924] = 18'b111111111111101101;
    mem[925] = 18'b111111111111110100;
    mem[926] = 18'b000000000000000100;
    mem[927] = 18'b111111111111110101;
    mem[928] = 18'b000000000000000101;
    mem[929] = 18'b000000000000000101;
    mem[930] = 18'b000000000000000001;
    mem[931] = 18'b000000000000000110;
    mem[932] = 18'b000000000000011100;
    mem[933] = 18'b111111111111111000;
    mem[934] = 18'b111111111111111001;
    mem[935] = 18'b000000000000010011;
    mem[936] = 18'b111111111111111011;
    mem[937] = 18'b111111111111101101;
    mem[938] = 18'b111111111111111111;
    mem[939] = 18'b000000000000000001;
    mem[940] = 18'b000000000000001001;
    mem[941] = 18'b000000000000000111;
    mem[942] = 18'b000000000000011111;
    mem[943] = 18'b000000000000001010;
    mem[944] = 18'b000000000000000011;
    mem[945] = 18'b111111111111101101;
    mem[946] = 18'b000000000000000111;
    mem[947] = 18'b000000000000010101;
    mem[948] = 18'b111111111111111000;
    mem[949] = 18'b000000000000010001;
    mem[950] = 18'b111111111111111011;
    mem[951] = 18'b000000000000011010;
    mem[952] = 18'b000000000000011001;
    mem[953] = 18'b000000000000001101;
    mem[954] = 18'b000000000000001000;
    mem[955] = 18'b000000000000011001;
    mem[956] = 18'b111111111111111101;
    mem[957] = 18'b000000000000001010;
    mem[958] = 18'b000000000000010000;
    mem[959] = 18'b000000000000000011;
    mem[960] = 18'b000000000000001110;
    mem[961] = 18'b000000000000010000;
    mem[962] = 18'b000000000000000101;
    mem[963] = 18'b000000000000000111;
    mem[964] = 18'b000000000000010000;
    mem[965] = 18'b000000000000010010;
    mem[966] = 18'b000000000000000101;
    mem[967] = 18'b000000000000000011;
    mem[968] = 18'b000000000000001011;
    mem[969] = 18'b000000000000000001;
    mem[970] = 18'b111111111111110000;
    mem[971] = 18'b111111111111110100;
    mem[972] = 18'b000000000000000101;
    mem[973] = 18'b000000000000001010;
    mem[974] = 18'b000000000000000010;
    mem[975] = 18'b000000000000010000;
    mem[976] = 18'b000000000000010011;
    mem[977] = 18'b111111111111110001;
    mem[978] = 18'b111111111111101111;
    mem[979] = 18'b000000000000011100;
    mem[980] = 18'b000000000000001010;
    mem[981] = 18'b000000000000000110;
    mem[982] = 18'b111111111111111011;
    mem[983] = 18'b000000000000010101;
    mem[984] = 18'b111111111111110011;
    mem[985] = 18'b000000000000000100;
    mem[986] = 18'b111111111111110100;
    mem[987] = 18'b000000000000001000;
    mem[988] = 18'b000000000000000001;
    mem[989] = 18'b111111111111111100;
    mem[990] = 18'b000000000000001101;
    mem[991] = 18'b000000000000000010;
    mem[992] = 18'b111111111111111111;
    mem[993] = 18'b000000000000000111;
    mem[994] = 18'b111111111111111100;
    mem[995] = 18'b000000000000010100;
    mem[996] = 18'b000000000000001010;
    mem[997] = 18'b000000000000000001;
    mem[998] = 18'b000000000000010010;
    mem[999] = 18'b000000000000000000;
    mem[1000] = 18'b000000000000010111;
    mem[1001] = 18'b000000000000000110;
    mem[1002] = 18'b000000000000010000;
    mem[1003] = 18'b111111111111111111;
    mem[1004] = 18'b111111111111111011;
    mem[1005] = 18'b111111111111111111;
    mem[1006] = 18'b111111111111101110;
    mem[1007] = 18'b111111111111011011;
    mem[1008] = 18'b000000000000101000;
    mem[1009] = 18'b000000000000010010;
    mem[1010] = 18'b111111111111100110;
    mem[1011] = 18'b000000000000011010;
    mem[1012] = 18'b000000000000010010;
    mem[1013] = 18'b000000000000001110;
    mem[1014] = 18'b000000000000111000;
    mem[1015] = 18'b000000000000001010;
    mem[1016] = 18'b000000000000101111;
    mem[1017] = 18'b111111111111111100;
    mem[1018] = 18'b111111111111111010;
    mem[1019] = 18'b111111111111111001;
    mem[1020] = 18'b000000000000011101;
    mem[1021] = 18'b000000000000011000;
    mem[1022] = 18'b000000000000011001;
    mem[1023] = 18'b000000000000001000;
    mem[1024] = 18'b111111111111101001;
    mem[1025] = 18'b000000000000010100;
    mem[1026] = 18'b111111111111111100;
    mem[1027] = 18'b111111111111110010;
    mem[1028] = 18'b111111111111110010;
    mem[1029] = 18'b000000000000000110;
    mem[1030] = 18'b000000000000001101;
    mem[1031] = 18'b000000000000000111;
    mem[1032] = 18'b111111111111101101;
    mem[1033] = 18'b111111111111110010;
    mem[1034] = 18'b000000000000010100;
    mem[1035] = 18'b111111111111101111;
    mem[1036] = 18'b111111111111110111;
    mem[1037] = 18'b000000000000000111;
    mem[1038] = 18'b000000000000100001;
    mem[1039] = 18'b000000000000011111;
    mem[1040] = 18'b000000000000000000;
    mem[1041] = 18'b111111111111111101;
    mem[1042] = 18'b000000000000000100;
    mem[1043] = 18'b111111111111101001;
    mem[1044] = 18'b111111111111100110;
    mem[1045] = 18'b111111111111101110;
    mem[1046] = 18'b111111111111101011;
    mem[1047] = 18'b000000000000011111;
    mem[1048] = 18'b000000000000000110;
    mem[1049] = 18'b111111111111010010;
    mem[1050] = 18'b000000000000000111;
    mem[1051] = 18'b111111111111111110;
    mem[1052] = 18'b111111111111100100;
    mem[1053] = 18'b111111111111101001;
    mem[1054] = 18'b000000000000010100;
    mem[1055] = 18'b000000000000001100;
    mem[1056] = 18'b000000000000100011;
    mem[1057] = 18'b000000000000010001;
    mem[1058] = 18'b000000000000000110;
    mem[1059] = 18'b111111111111101010;
    mem[1060] = 18'b000000000000010111;
    mem[1061] = 18'b000000000000000001;
    mem[1062] = 18'b111111111111110011;
    mem[1063] = 18'b000000000000010010;
    mem[1064] = 18'b000000000000000100;
    mem[1065] = 18'b000000000000000101;
    mem[1066] = 18'b000000000000001110;
    mem[1067] = 18'b000000000000011000;
    mem[1068] = 18'b111111111111111111;
    mem[1069] = 18'b000000000000010111;
    mem[1070] = 18'b000000000000101010;
    mem[1071] = 18'b000000000000001110;
    mem[1072] = 18'b000000000000010111;
    mem[1073] = 18'b000000000000001100;
    mem[1074] = 18'b000000000000010001;
    mem[1075] = 18'b000000000000000011;
    mem[1076] = 18'b000000000000001011;
    mem[1077] = 18'b000000000000011000;
    mem[1078] = 18'b000000000000001000;
    mem[1079] = 18'b111111111111111110;
    mem[1080] = 18'b111111111111111011;
    mem[1081] = 18'b000000000000001001;
    mem[1082] = 18'b000000000000010111;
    mem[1083] = 18'b000000000000101110;
    mem[1084] = 18'b000000000000001010;
    mem[1085] = 18'b000000000000000111;
    mem[1086] = 18'b000000000000010100;
    mem[1087] = 18'b000000000000001010;
    mem[1088] = 18'b000000000000000111;
    mem[1089] = 18'b000000000000011111;
    mem[1090] = 18'b000000000000001010;
    mem[1091] = 18'b000000000001110100;
    mem[1092] = 18'b000000000000000101;
    mem[1093] = 18'b000000000000001011;
    mem[1094] = 18'b000000000000000000;
    mem[1095] = 18'b000000000000100001;
    mem[1096] = 18'b000000000000000100;
    mem[1097] = 18'b111111111111111111;
    mem[1098] = 18'b000000000000000010;
    mem[1099] = 18'b111111111111110000;
    mem[1100] = 18'b111111111111011111;
    mem[1101] = 18'b111111111111111011;
    mem[1102] = 18'b000000000000001010;
    mem[1103] = 18'b000000000000001110;
    mem[1104] = 18'b111111111111111001;
    mem[1105] = 18'b111111111111011011;
    mem[1106] = 18'b111111111111110100;
    mem[1107] = 18'b111111111111111101;
    mem[1108] = 18'b111111111111110110;
    mem[1109] = 18'b000000000000001001;
    mem[1110] = 18'b000000000000000010;
    mem[1111] = 18'b000000000000000101;
    mem[1112] = 18'b000000000000010101;
    mem[1113] = 18'b000000000000001011;
    mem[1114] = 18'b000000000000000011;
    mem[1115] = 18'b000000000000011000;
    mem[1116] = 18'b000000000000000100;
    mem[1117] = 18'b000000000000010000;
    mem[1118] = 18'b000000000000000101;
    mem[1119] = 18'b000000000000000000;
    mem[1120] = 18'b111111111111111110;
    mem[1121] = 18'b000000000000001010;
    mem[1122] = 18'b000000000000000010;
    mem[1123] = 18'b000000000000001010;
    mem[1124] = 18'b000000000000000110;
    mem[1125] = 18'b111111111111111110;
    mem[1126] = 18'b000000000000001010;
    mem[1127] = 18'b000000000000001010;
    mem[1128] = 18'b111111111111110011;
    mem[1129] = 18'b000000000000001101;
    mem[1130] = 18'b000000000000001000;
    mem[1131] = 18'b111111111111110010;
    mem[1132] = 18'b111111111111101111;
    mem[1133] = 18'b111111111111111010;
    mem[1134] = 18'b111111111111101011;
    mem[1135] = 18'b000000000000000010;
    mem[1136] = 18'b000000000000010000;
    mem[1137] = 18'b000000000000010000;
    mem[1138] = 18'b000000000000001011;
    mem[1139] = 18'b000000000000000001;
    mem[1140] = 18'b000000000000010011;
    mem[1141] = 18'b111111111111110101;
    mem[1142] = 18'b000000000000101000;
    mem[1143] = 18'b111111111111100101;
    mem[1144] = 18'b111111111111111011;
    mem[1145] = 18'b111111111111110110;
    mem[1146] = 18'b111111111111101110;
    mem[1147] = 18'b111111111111111111;
    mem[1148] = 18'b111111111111100010;
    mem[1149] = 18'b111111111111110000;
    mem[1150] = 18'b000000000000001001;
    mem[1151] = 18'b111111111111111011;
    mem[1152] = 18'b111111111111111011;
    mem[1153] = 18'b111111111111111101;
    mem[1154] = 18'b000000000000000110;
    mem[1155] = 18'b111111111111101010;
    mem[1156] = 18'b111111111111101101;
    mem[1157] = 18'b000000000101011000;
    mem[1158] = 18'b000000000100111011;
    mem[1159] = 18'b000000000100111010;
    mem[1160] = 18'b000000000010011001;
    mem[1161] = 18'b000000000000010011;
    mem[1162] = 18'b111111111111011010;
    mem[1163] = 18'b000000000000001001;
    mem[1164] = 18'b111111111111111110;
    mem[1165] = 18'b000000000000000100;
    mem[1166] = 18'b000000000000000010;
    mem[1167] = 18'b000000000000000001;
    mem[1168] = 18'b111111111111111011;
    mem[1169] = 18'b000000000000000010;
    mem[1170] = 18'b000000000000000100;
    mem[1171] = 18'b000000000000000011;
    mem[1172] = 18'b111111111111111110;
    mem[1173] = 18'b000000000000000100;
    mem[1174] = 18'b111111111111110111;
    mem[1175] = 18'b111111111111111011;
    mem[1176] = 18'b111111111111111110;
    mem[1177] = 18'b000000000000001010;
    mem[1178] = 18'b000000000000000010;
    mem[1179] = 18'b111111111111111011;
    mem[1180] = 18'b000000000000000100;
    mem[1181] = 18'b000000000000000111;
    mem[1182] = 18'b111111111111111001;
    mem[1183] = 18'b111111111111111110;
    mem[1184] = 18'b111111111111111000;
    mem[1185] = 18'b000000000000000011;
    mem[1186] = 18'b000000000000000011;
    mem[1187] = 18'b111111111111111010;
    mem[1188] = 18'b111111111111111000;
    mem[1189] = 18'b111111111111100110;
    mem[1190] = 18'b111111111111101010;
    mem[1191] = 18'b111111111111111001;
    mem[1192] = 18'b000000000000000001;
    mem[1193] = 18'b000000000000000011;
    mem[1194] = 18'b000000000000011110;
    mem[1195] = 18'b000000000000011111;
    mem[1196] = 18'b000000000000110111;
    mem[1197] = 18'b111111111111011100;
    mem[1198] = 18'b000000000011101010;
    mem[1199] = 18'b111111111111011110;
    mem[1200] = 18'b111111111111111101;
    mem[1201] = 18'b000000000000001110;
    mem[1202] = 18'b000000000000001010;
    mem[1203] = 18'b111111111111111101;
    mem[1204] = 18'b000000000000001000;
    mem[1205] = 18'b000000000000000100;
    mem[1206] = 18'b111111111111111110;
    mem[1207] = 18'b000000000000000110;
    mem[1208] = 18'b111111111111110110;
    mem[1209] = 18'b000000000000001001;
    mem[1210] = 18'b111111111111111101;
    mem[1211] = 18'b000000000000001100;
    mem[1212] = 18'b000000000100100011;
    mem[1213] = 18'b000000000100111000;
    mem[1214] = 18'b000000000101011010;
    mem[1215] = 18'b000000000011000101;
    mem[1216] = 18'b111111111111010100;
    mem[1217] = 18'b000000000001111010;
    mem[1218] = 18'b111111111111110010;
    mem[1219] = 18'b000000000000000010;
    mem[1220] = 18'b111111111111111011;
    mem[1221] = 18'b000000000001000010;
    mem[1222] = 18'b000000000000100000;
    mem[1223] = 18'b000000000000001010;
    mem[1224] = 18'b000000000000000110;
    mem[1225] = 18'b000000000000000110;
    mem[1226] = 18'b000000000000001101;
    mem[1227] = 18'b000000000000000001;
    mem[1228] = 18'b000000000000000101;
    mem[1229] = 18'b000000000000001000;
    mem[1230] = 18'b000000000000000100;
    mem[1231] = 18'b000000000000000001;
    mem[1232] = 18'b111111111111110101;
    mem[1233] = 18'b000000000000000010;
    mem[1234] = 18'b000000000000000101;
    mem[1235] = 18'b111111111111111110;
    mem[1236] = 18'b111111111111111001;
    mem[1237] = 18'b000000000000000010;
    mem[1238] = 18'b000000000000000001;
    mem[1239] = 18'b111111111111111111;
    mem[1240] = 18'b000000000000001100;
    mem[1241] = 18'b111111111111111010;
    mem[1242] = 18'b111111111111111010;
    mem[1243] = 18'b000000000000000011;
    mem[1244] = 18'b000000000000001001;
    mem[1245] = 18'b000000000000000110;
    mem[1246] = 18'b000000000000000010;
    mem[1247] = 18'b000000000000001001;
    mem[1248] = 18'b111111111111111111;
    mem[1249] = 18'b000000000000000100;
    mem[1250] = 18'b000000000000000000;
    mem[1251] = 18'b111111111111111100;
    mem[1252] = 18'b111111111111111011;
    mem[1253] = 18'b111111111111111110;
    mem[1254] = 18'b000000000000000010;
    mem[1255] = 18'b111111111111111010;
    mem[1256] = 18'b000000000000000100;
    mem[1257] = 18'b000000000000001101;
    mem[1258] = 18'b000000000000000000;
    mem[1259] = 18'b111111111111111100;
    mem[1260] = 18'b111111111100001101;
    mem[1261] = 18'b111111111111110011;
    mem[1262] = 18'b000000000001010001;
    mem[1263] = 18'b111111111111110010;
    mem[1264] = 18'b111111111111110110;
    mem[1265] = 18'b000000000000000100;
    mem[1266] = 18'b000000000010011001;
    mem[1267] = 18'b000000000011000010;
    mem[1268] = 18'b000000000001111101;
    mem[1269] = 18'b111111111111111010;
    mem[1270] = 18'b000000000100111011;
    mem[1271] = 18'b000000000011011111;
    mem[1272] = 18'b111111111111111001;
    mem[1273] = 18'b111111111111111110;
    mem[1274] = 18'b111111111111111111;
    mem[1275] = 18'b000000000000000000;
    mem[1276] = 18'b111111111111111110;
    mem[1277] = 18'b000000000000000010;
    mem[1278] = 18'b000000000000000010;
    mem[1279] = 18'b111111111111111111;
    mem[1280] = 18'b111111111111111000;
    mem[1281] = 18'b111111111111111001;
    mem[1282] = 18'b111111111111111111;
    mem[1283] = 18'b111111111111111011;
    mem[1284] = 18'b000000000011100111;
    mem[1285] = 18'b000000000011010110;
    mem[1286] = 18'b000000000011000001;
    mem[1287] = 18'b000000000011110011;
    mem[1288] = 18'b000000000000001010;
    mem[1289] = 18'b111111111111111010;
    mem[1290] = 18'b000000000000100001;
    mem[1291] = 18'b111111111111011001;
    mem[1292] = 18'b000000000000101110;
    mem[1293] = 18'b000000000000001110;
    mem[1294] = 18'b000000000000010110;
    mem[1295] = 18'b111111111111110010;
    mem[1296] = 18'b111111111111111110;
    mem[1297] = 18'b111111111111110010;
    mem[1298] = 18'b000000000000000011;
    mem[1299] = 18'b111111111111111011;
    mem[1300] = 18'b111111111111111100;
    mem[1301] = 18'b111111111111111000;
    mem[1302] = 18'b000000000000000010;
    mem[1303] = 18'b000000000000000001;
    mem[1304] = 18'b000000000000000000;
    mem[1305] = 18'b000000000000001000;
    mem[1306] = 18'b000000000000000001;
    mem[1307] = 18'b000000000000000000;
    mem[1308] = 18'b111111111111111111;
    mem[1309] = 18'b111111111111111001;
    mem[1310] = 18'b000000000000001011;
    mem[1311] = 18'b000000000000000100;
    mem[1312] = 18'b111111111111111111;
    mem[1313] = 18'b111111111111111100;
    mem[1314] = 18'b000000000000000000;
    mem[1315] = 18'b000000000000000011;
    mem[1316] = 18'b111111111111111010;
    mem[1317] = 18'b000000000000000001;
    mem[1318] = 18'b000000000000000010;
    mem[1319] = 18'b000000000000000001;
    mem[1320] = 18'b000000000000000101;
    mem[1321] = 18'b000000000000000010;
    mem[1322] = 18'b111111111111111101;
    mem[1323] = 18'b111111111111111100;
    mem[1324] = 18'b111111111111111101;
    mem[1325] = 18'b000000000000000000;
    mem[1326] = 18'b111111111111111100;
    mem[1327] = 18'b111111111111111110;
    mem[1328] = 18'b000000000000000001;
    mem[1329] = 18'b000000000000000010;
    mem[1330] = 18'b000000000000001011;
    mem[1331] = 18'b000000000000000011;
    mem[1332] = 18'b000000000000000001;
    mem[1333] = 18'b000000000000000011;
    mem[1334] = 18'b000000000000000110;
    mem[1335] = 18'b000000000000000001;
    mem[1336] = 18'b111111111111111101;
    mem[1337] = 18'b000000000000000101;
    mem[1338] = 18'b111111111111111111;
    mem[1339] = 18'b111111111111110101;
    mem[1340] = 18'b000000000000000101;
    mem[1341] = 18'b000000000000001000;
    mem[1342] = 18'b111111111111111100;
    mem[1343] = 18'b111111111111111110;
    mem[1344] = 18'b000000000000000000;
    mem[1345] = 18'b000000000000000000;
    mem[1346] = 18'b000000000000000000;
    mem[1347] = 18'b000000000000000000;
    mem[1348] = 18'b000000000000000000;
    mem[1349] = 18'b000000000000000000;
    mem[1350] = 18'b000000000000000000;
    mem[1351] = 18'b000000000000000000;
    mem[1352] = 18'b000000000000000000;
    mem[1353] = 18'b000000000000000000;
    mem[1354] = 18'b000000000000000000;
    mem[1355] = 18'b000000000000000000;
    mem[1356] = 18'b000000000000000000;
    mem[1357] = 18'b000000000000000000;
    mem[1358] = 18'b000000000000000000;
    mem[1359] = 18'b000000000000000000;
    mem[1360] = 18'b000000000000000000;
    mem[1361] = 18'b000000000000000000;
    mem[1362] = 18'b000000000000000000;
    mem[1363] = 18'b000000000000000000;
    mem[1364] = 18'b000000000000000000;
    mem[1365] = 18'b000000000000000000;
    mem[1366] = 18'b000000000000000000;
    mem[1367] = 18'b000000000000000000;
    mem[1368] = 18'b000000000000000000;
    mem[1369] = 18'b000000000000000000;
    mem[1370] = 18'b000000000000000000;
    mem[1371] = 18'b000000000000000000;
    mem[1372] = 18'b000000000000000000;
    mem[1373] = 18'b000000000000000000;
    mem[1374] = 18'b000000000000000000;
    mem[1375] = 18'b000000000000000000;
    mem[1376] = 18'b000000000000000000;
    mem[1377] = 18'b000000000000000000;
    mem[1378] = 18'b000000000000000000;
    mem[1379] = 18'b000000000000000000;
    mem[1380] = 18'b000000000000000000;
    mem[1381] = 18'b000000000000000000;
    mem[1382] = 18'b000000000000000000;
    mem[1383] = 18'b000000000000000000;
    mem[1384] = 18'b000000000000000000;
    mem[1385] = 18'b000000000000000000;
    mem[1386] = 18'b000000000000000000;
    mem[1387] = 18'b000000000000000000;
    mem[1388] = 18'b000000000000000000;
    mem[1389] = 18'b000000000000000000;
    mem[1390] = 18'b000000000000000000;
    mem[1391] = 18'b000000000000000000;
    mem[1392] = 18'b000000000000000000;
    mem[1393] = 18'b000000000000000000;
    mem[1394] = 18'b000000000000000000;
    mem[1395] = 18'b000000000000000000;
    mem[1396] = 18'b000000000000000000;
    mem[1397] = 18'b000000000000000000;
    mem[1398] = 18'b000000000000000000;
    mem[1399] = 18'b000000000000000000;
    mem[1400] = 18'b000000000000000000;
    mem[1401] = 18'b000000000000000000;
    mem[1402] = 18'b000000000000000000;
    mem[1403] = 18'b000000000000000000;
    mem[1404] = 18'b000000000000000000;
    mem[1405] = 18'b000000000000000000;
    mem[1406] = 18'b000000000000000000;
    mem[1407] = 18'b000000000000000000;
    mem[1408] = 18'b000000000000000000;
    mem[1409] = 18'b000000000000000000;
    mem[1410] = 18'b000000000000000000;
    mem[1411] = 18'b000000000000000000;
    mem[1412] = 18'b000000000000000000;
    mem[1413] = 18'b000000000000000000;
    mem[1414] = 18'b000000000000000000;
    mem[1415] = 18'b000000000000000000;
    mem[1416] = 18'b000000000000000000;
    mem[1417] = 18'b000000000000000000;
    mem[1418] = 18'b000000000000000000;
    mem[1419] = 18'b000000000000000000;
    mem[1420] = 18'b000000000000000000;
    mem[1421] = 18'b000000000000000000;
    mem[1422] = 18'b000000000000000000;
    mem[1423] = 18'b000000000000000000;
    mem[1424] = 18'b000000000000000000;
    mem[1425] = 18'b000000000000000000;
    mem[1426] = 18'b000000000000000000;
    mem[1427] = 18'b000000000000000000;
    mem[1428] = 18'b000000000000000000;
    mem[1429] = 18'b000000000000000000;
    mem[1430] = 18'b000000000000000000;
    mem[1431] = 18'b000000000000000000;
    mem[1432] = 18'b000000000000000000;
    mem[1433] = 18'b000000000000000000;
    mem[1434] = 18'b000000000000000000;
    mem[1435] = 18'b000000000000000000;
    mem[1436] = 18'b000000000000000000;
    mem[1437] = 18'b000000000000000000;
    mem[1438] = 18'b000000000000000000;
    mem[1439] = 18'b000000000000000000;
  end
  
endmodule