`include "num_data.v"

module w_rom_17 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b111111110110101111000000000110000111000000000101011001111111111001011111000000000000010110111111111110000111000000000100101111111111111010101011111111111000010110;
    mem[1] = 162'b111111110101000010111111110010000110000000000101110000000000000000111111000000000001110011111111111110110111111111110110110100000000000010100110111111111101101000;
    mem[2] = 162'b111111111101110001111111111110101011111111111101000110000000001001111100000000000110011010000000000001010110111111111000111001111111111010001001111111111001011000;
    mem[3] = 162'b111111110111001010000000000101101010000000000100011000111111111110011010000000000000101111000000000110000010111111110110100000111111111010011100000000000101000001;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111000111100111111111010110001000000000000101100000000000001000011111111111010100000111111111111001010111111111101110101111111111010101101000000000110100110;
    mem[33] = 162'b000000000110111010000000000000010100111111111111111110111111111100010010000000000001111110111111111010101011111111111111111101111111111001110101000000000000111000;
    mem[34] = 162'b111111110111101001111111111011010011111111110110110011000000000011111101111111111101001100111111111010000101111111111110101001111111111100111000111111111111100111;
    mem[35] = 162'b111111111100010101111111111100010011000000000010111010111111111100001001111111110111010100000000000001011110111111111011000111000000000100100011111111110111000011;
    mem[36] = 162'b111111111011010110111111111110011110000000000001010001000000000010101101000000000100101011000000000100001100000000000100100001111111111011100101000000000110000000;
    mem[37] = 162'b000000000000011011000000000001011101000000000010110101111111111000011001111111111001011101000000000111101110000000000000101100111111111101011000111111111011110001;
    mem[38] = 162'b000000000111001111000000001000001001111111111110011010111111111110001010000000000001001001000000000101111111000000000101000011000000000001100111000000000111110000;
    mem[39] = 162'b111111111001000010000000000100000000000000001000101000111111111101001001000000000000001000111111111101101111111111111101111000000000000110101100111111111011111011;
    mem[40] = 162'b111111111001010101000000000111100101000000000100001011000000001000101110000000000011011000000000000101101110000000000001001111000000000000110111000000000011101111;
    mem[41] = 162'b000000000110010000000000000001111010111111111100001101111111111010110100000000000000110100000000000001100011111111111101011110000000000111111001000000000010011010;
    mem[42] = 162'b000000000100000011000000000001100110111111111100001000000000000001011111000000000011100011000000000000000010000000000000010101111111101111111110000000000110101001;
    mem[43] = 162'b111111111001001110000000000010010111111111111010011000111111111010101111000000000010011010000000000010110010000000000110011001111111111101001000000000000101100110;
    mem[44] = 162'b111111111110101101111111111101001100000000000100101010000000000110010110000000000000000101111111111100011001111111111100001110000000000111100111000000000000000111;
    mem[45] = 162'b000000000101010001000000000010001001111111111101010001000000000010101010000000000011000000111111111111010010111111111011010001111111111100011010111111111111100000;
    mem[46] = 162'b000000000110011011000000001011001011000000000101100011000000000011110110111111111000110001111111111010100111111111110011110101000000000010110010111111111111010100;
    mem[47] = 162'b000000000011000011000000001000111001111111111101101000111111111011101011111111111110011100111111111011011011000000000001001111000000000011110101111111111111101100;
    mem[48] = 162'b000000000011111101111111111100000100000000000011101100000000000000011111111111111010100101111111111111101001111111111111111110000000000010000101000000000000101011;
    mem[49] = 162'b000000000011000001111111111110110001111111111001110100000000000000100010111111111101000001000000000101110010111111111110011010111111111110111100111111110110001001;
    mem[50] = 162'b000000000000111010111111111001110010111111111110010011111111110011110010000000000001100110000000000000010011111111111011010110111111110110100100000000001111111100;
    mem[51] = 162'b000000000110111100000000000101010011111111111110001100000000001010110111000000000001000001000000000110111000000000000100100100000000001000010101000000000011101010;
    mem[52] = 162'b000000000011101100111111111110011011000000000110101100000000000110110110000000000001010001111111111100101000000000001000011001000000000110011011111111111011010000;
    mem[53] = 162'b111111111111010000000000000000000110000000000010001100111111111110000010111111111101011101111111110011010001000000000110101100000000000101000111111111111101101101;
    mem[54] = 162'b111111111110000100111111111011001110000000000011001111111111111110100111111111111110110110111111111111101000000000000011011100000000000011101001000000000011001111;
    mem[55] = 162'b111111111111000010111111111111101001111111110101010100111111111000000001000000000010101101000000000001011101000000000001111111111111111001110100000000000100011100;
    mem[56] = 162'b000000000001111110111111111100111101000000000001011011111111111111110001000000000000001101111111111010110100111111111000100011000000000011100010111111111111101010;
    mem[57] = 162'b000000000001110011000000000000101110111111111010011001000000000000011101000000000101110010000000000010011101000000001001101111111111110011010110111111111010111100;
    mem[58] = 162'b111111111010111111111111111100101111111111111110101001111111111001101101111111111011011010111111111101101101000000001001010010111111111111100101000000000000111110;
    mem[59] = 162'b000000000101000011111111111110010000111111111010001110000000000000011101111111111111011001111111111110011011000000000111101111111111111001101001111111110100100000;
    mem[60] = 162'b000000000011100010000000000010001001000000000011101100000000000011101101000000000010011001000000000100000010000000000010001101111111110111001010111111110101110110;
    mem[61] = 162'b000000000010000111111111111100100100111111111111100111111111111111010010111111111110110010000000000110110001000000000100110100000000000101111111111111111011111110;
    mem[62] = 162'b111111111101001110111111111110010000000000001000100000000000000111010110000000000010010111000000000000000100111111111011000100000000000001010011111111110101101100;
    mem[63] = 162'b000000000110110111000000000100000110111111111110111101111111111100011011111111111110101110000000000010101010000000000011101101000000000010110000000000000011111010;
    mem[64] = 162'b000000000011001011000000000110001101111111111011011111111111111111100011111111111111011010000000000011011100000000000110001010111111111010100100111111110010001010;
    mem[65] = 162'b111111111100011101000000000000100001111111111100100011000000000010010111111111111001011101000000000000101001000000001011010100000000000101110100000000000100000011;
    mem[66] = 162'b111111111010011101111111111110111101111111111011010011000000000011000001000000000010101011111111111111010100000000000000011100000000000010100000111111111011100111;
    mem[67] = 162'b111111111100100010111111111101010011111111111111001010000000000101000010111111111001101111000000000001010011111111111101101011000000000001110011000000000001101111;
    mem[68] = 162'b111111111110000101111111111101111000000000000000100110111111111110000010111111111001111011000000000000110000000000000000100011000000000001001000111111111101110001;
    mem[69] = 162'b111111111010111101000000000011000111000000000010111010000000000100001011111111111100111110000000000000110101000000000010101100000000000101100111000000000010010001;
    mem[70] = 162'b000000000010110011000000000000111100111111111110101110000000000100010110111111111011110110000000000101001011000000000010101010000000000000111001000000000000000010;
    mem[71] = 162'b000000000001000011111111111100001100000000000000010010000000001010000100000000000000011110111111111111001000000000000010001111111111111110000110000000000001011010;
    mem[72] = 162'b111111111010101011111111111110111010111111111010011010000000000010110001111111111100101000111111111101000101000000000011111101111111111111011010111111111110111001;
    mem[73] = 162'b000000000000100101111111111010100111111111111111101010000000000011001011111111111011001010111111111111100101000000000111001110111111111100110000000000000000111101;
    mem[74] = 162'b111111111111000001000000000011101110000000000100101010000000000011000010111111111111100001111111111111010100111111111001010101111111111111110001000000000010001101;
    mem[75] = 162'b000000000011110101000000000000011111000000000100010011000000000000011110000000000001100011000000000010010111111111111110001101000000000000010001111111111101001111;
    mem[76] = 162'b000000000110100011000000000111010111000000000001011111000000000000100010000000000111110000111111111111010010000000000100101000000000000011000010000000000010101000;
    mem[77] = 162'b000000000010100000111111111101010101000000000010110001111111111101101001111111111110110001111111111011100100000000000001101100000000000000000101000000000000001101;
    mem[78] = 162'b000000001001001011000000000100001111000000000010000101000000001010010010000000000111001110000000000011011011000000000100010001000000000110000001111111111100001100;
    mem[79] = 162'b111111111101000101111111111110010100000000000000011101111111111001001110000000000011100000111111111100101110111111111111110000111111111011111101111111111010111101;
    mem[80] = 162'b111111111000001010111111111010100100111111111110100011111111111100010111111111111011010010000000000001010011000000000010110100111111111011010110111111111101111111;
    mem[81] = 162'b111111111110011110111111111001100001111111111111011100111111111000101100000000000010100000111111111111001100000000000011111010111111111010111010111111111110100110;
    mem[82] = 162'b000000000011111001000000000110001000111111111111000001000000000101000000111111111110000011111111111100111100000000000101010110000000000001111100111111111111100011;
    mem[83] = 162'b000000000001011011000000000001100000000000000100011110000000000001010100000000000001110100111111111011100100000000000001110011000000000110001011111111111100001010;
    mem[84] = 162'b111111111111100000111111111111000011111111111111101100000000000010010100111111111100010011111111111100001001111111111011001101111111111101110111111111111110101100;
    mem[85] = 162'b000000001000101001000000000000101000111111111010001110000000001001110111000000000001100100000000000100111001000000000001011100000000000001001000000000000000100101;
    mem[86] = 162'b000000000000010110000000000001110010000000000100100001000000001001001000000000000011011110000000000101000010000000000111000100000000000110010100000000000010001100;
    mem[87] = 162'b000000000000110111000000000000111001111111111111111100111111111110101111000000000000001000111111111011101111111111111001100100111111111010001101111111110111011110;
    mem[88] = 162'b000000000001011110111111111111111001111111111001110001000000000001011010111111111110110110000000000000100001000000000001001110000000000011000100111111111001100011;
    mem[89] = 162'b111111111101010110111111111100001010111111111011010111111111111100100101000000000011010011000000000001101001000000000000010011111111111111101001000000000100110011;
    mem[90] = 162'b111111111100000110000000000011001101111111111110001010111111111110010001000000000001000000111111111111101100000000000000000100000000000100000100000000000001010111;
    mem[91] = 162'b111111111111111010000000000001111111000000000011110101000000000110001011111111111011100011111111111001101101000000000100100000111111111011100001111111111101010100;
    mem[92] = 162'b000000000001100011111111111100001111111111111101111111111111110111001010111111111111011000000000000011000000000000000000011011111111111101101100000000000010110001;
    mem[93] = 162'b000000000000101011111111111110000111111111111011110011111111111100111011000000000000100001000000000101100011111111110110111001000000000010000110111111111110111101;
    mem[94] = 162'b111111111101110111111111111101000001000000000010110101111111111101000100000000000001111100111111111011110111000000000000100100111111111101010001000000000101110000;
    mem[95] = 162'b111111111111110100000000000000000001000000000011010000000000000001011100000000000000001000111111111110011000000000000011111010111111111101100000111111111100111101;
    mem[96] = 162'b111111111111111000111111111111111010000000000000010010000000000000000111111111111111111101111111111111101100111111111111111001111111111111111010000000000000010010;
    mem[97] = 162'b000000000000010001111111111111110010111111111111101111000000000000010100111111111111111110000000000000001101111111111111111001111111111111110001000000000000001110;
    mem[98] = 162'b111111111111011110000000000000001001111111111111111000000000000000001111000000000000011011000000000000001000111111111111101000111111111111110100111111111111111010;
    mem[99] = 162'b000000000000001100000000000000010000111111111111111011111111111111110111111111111111110111111111111111110001111111111111110111111111111111110000111111111111110111;
    mem[100] = 162'b111111111111101110111111111111111001111111111111101110111111111111111101000000000000000011111111111111111001000000000000000011111111111111111111111111111111111100;
    mem[101] = 162'b111111111111111111000000000000000001000000000000011010111111111111110011111111111111101101111111111111111010111111111111111000111111111111111100000000000000001001;
    mem[102] = 162'b000000000000001000000000000000010110000000000000010011111111111111111110000000000000001001111111111111111111111111111111111101111111111111110111000000000000000100;
    mem[103] = 162'b111111111111111000000000000000001011000000000000000111111111111111110111000000000000010001000000000000000000000000000000001110000000000000001100000000000000001001;
    mem[104] = 162'b111111111111111001111111111111110110111111111111111010000000000000001001111111111111101011111111111111110110000000000000000111111111111111110101000000000000000011;
    mem[105] = 162'b000000000000001010111111111111101111000000000000000100111111111111111110000000000000000010111111111111110101000000000000100010111111111111111010000000000000001101;
    mem[106] = 162'b000000000000000110000000000000001101000000000000000100111111111111111110000000000000000010000000000000000000000000000000000000111111111111111101000000000000000001;
    mem[107] = 162'b000000000000000001111111111111111001000000000000000110000000000000000011000000000000000111000000000000001110000000000000001100000000000000000010111111111111111011;
    mem[108] = 162'b111111111111111011111111111111110001111111111111110101111111111111111001000000000000000010111111111111110011000000000000000011111111111111110111111111111111111010;
    mem[109] = 162'b000000000000010100000000000000011000000000000000000001111111111111110111111111111111111100000000000000001010000000000000000010111111111111111001111111111111110011;
    mem[110] = 162'b000000000000000000000000000000001111111111111111111001111111111111111100000000000000000110111111111111110111000000000000000000000000000000000101111111111111111000;
    mem[111] = 162'b000000000000001100000000000000001000000000000000011101111111111111110110111111111111111001111111111111110110111111111111111101000000000000000010000000000000001000;
    mem[112] = 162'b000000000000101010000000000000010101111111111111101110000000000000001001000000000000000010000000000000001011000000000001011100000000000000010101111111111111111110;
    mem[113] = 162'b000000000000001110111111111111111100000000000000010101000000000000001110000000000000000000000000000000000011000000000000000011000000000000001000000000000000000000;
    mem[114] = 162'b000000000000001100000000000000001100111111111111111001000000000000000111000000000000001001000000000000001100000000000000001111000000000000000011111111111111110111;
    mem[115] = 162'b111111111111111100111111111111110101000000000000000010111111111111111011000000000000000010000000000000000100000000000000000100111111111111111000000000000000001010;
    mem[116] = 162'b000000000000000010111111111111111010000000000000000001111111111111111100111111111111110111111111111111111011111111111111111000111111111111110000111111111111111010;
    mem[117] = 162'b111111111111110110111111111111101010111111111111101000000000000000010010000000000000000011111111111111111001111111111111110111111111111111111000111111111111101100;
    mem[118] = 162'b111111111111111010111111111111111010111111111111111001111111111111111010111111111111100011111111111111110011111111111111111111111111111111111110000000000000001110;
    mem[119] = 162'b000000000000000110000000000000001000000000000000001001000000000000000000000000000000000000000000000000001000000000000000000011111111111111101100000000000000001101;
    mem[120] = 162'b000000000000000101111111111111110001000000000000010001000000000000001111111111111111111111000000000000010000111111111111111101111111111111101111111111111111111011;
    mem[121] = 162'b000000000000001111111111111111111111000000000000100011000000000000000100111111111111111110000000000000001100111111111111010111111111111111101100000000000000000101;
    mem[122] = 162'b000000000000010101000000000000000001111111111111111010000000000000000000111111111111110000111111111111111101000000000000010001000000000000001100000000000000001100;
    mem[123] = 162'b111111111111111001111111111111111011000000000000000011111111111111110010111111111111111001111111111111111010111111111111111000111111111111111100111111111111111011;
    mem[124] = 162'b000000000000001011000000000000000010111111111111111001111111111111111110111111111111111011111111111111111100111111111111110110111111111111101010111111111111101010;
    mem[125] = 162'b111111111111111000111111111111111110111111111111101101000000000000001100000000000000000110000000000000001001000000000000000001000000000000000000111111111111111100;
    mem[126] = 162'b000000000000000101111111111111110001111111111111110101000000000000000101111111111111111011000000000000010000000000000000000110000000000000011110000000000000001110;
    mem[127] = 162'b111111111111110110000000000000000011111111111111111110000000000000000010000000000000001000111111111111110101111111111111111011000000000000000000111111111111111101;
    mem[128] = 162'b000000000000011001000000000101000111000000000101000111000000000100101000000000000000110011000000000000010110000000000000000010000000000000100101111111111111110100;
    mem[129] = 162'b000000000000000100000000000000001100000000000000000100111111111111110110000000000000000010000000000000001100000000000001111011111111111111110000111111111111010010;
    mem[130] = 162'b000000000000000110000000000000000011111111111111111010000000000000001010111111111111111010000000000000000111000000000000001000111111111111111101111111111111111101;
    mem[131] = 162'b111111111111111110111111111111111110000000000000000110000000000000000100000000000000001101000000000000000010000000000000000100000000000000001000000000000000001011;
    mem[132] = 162'b111111111111111101111111111111100110000000000000100001000000000000000001000000000000001110111111111111110110111111111111101101111111111111110110000000000000001110;
    mem[133] = 162'b111111111111111111000000000000001011000000000000000100000000000000000100000000000000000111000000000000001001111111111111100100111111111111110101111111111111101001;
    mem[134] = 162'b000000000010110110000000000101110101000000000100101011000000000000001100000000000000000001000000000000001110000000000000001001000000000000001000111111111111111001;
    mem[135] = 162'b000000000001000101111111111111111100111111111111110100000000000000010100000000000000000000000000000001101111111111111111111110000000000000010001000000000100011110;
    mem[136] = 162'b000000000000001100111111111111111111111111111111111101111111111111111011000000000000000101000000000000000011111111111111111101111111111111111111000000000000000111;
    mem[137] = 162'b000000000000001100000000000000010101111111111111111011000000000000010000000000000000010010000000000000001000000000000000001100000000000000001111000000000000000111;
    mem[138] = 162'b000000000000000100111111111111111110000000000000000001000000000000000100000000000000001000000000000000011001000000000000001110000000000000010101000000000000001111;
    mem[139] = 162'b000000000000000100111111111111111111000000000000001111000000000000000111000000000000000100000000000000001011000000000000000101000000000000000111000000000000000101;
    mem[140] = 162'b000000000010011000000000000100101000000000000101011001000000000001111111000000000000111110111111111111100001111111111111011010000000000000010000111111111101100001;
    mem[141] = 162'b111111111111110110111111111111111001111111111111111110111111111111110001000000000000001010000000000000000101000000000100010011000000000001000101000000000011010111;
    mem[142] = 162'b000000000100100111000000000100110111000000000010110101111111111111110010111111111111110100111111111111111001111111111111101111000000000000000101111111111111110010;
    mem[143] = 162'b000000000000110110111111111111101100111111111111011011000000000000001010111111111111110000111111111111111110111111111111011010000000000000010110000000000010001111;
    mem[144] = 162'b111111111111111011111111111111111011111111111111110001111111111111111010111111111111101101111111111111111010111111111111111011111111111111110111000000000000000000;
    mem[145] = 162'b111111111111111011000000000000000011111111111111110111111111111111111001000000000000000011000000000000000010111111111111111001111111111111111001000000000000000011;
    mem[146] = 162'b000000000000000001111111111111111010111111111111110110000000000000000000111111111111111010000000000000000101000000000000000001000000000000000110111111111111111000;
    mem[147] = 162'b000000000000000011000000000000000100000000000000010001000000000000000000000000000000000110000000000000000001111111111111111111000000000000000000000000000000001111;
    mem[148] = 162'b000000000000000100000000000000001000000000000000000100000000000000000110000000000000000011000000000000011100000000000000001001000000000000000100000000000000001101;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111101000000000000001001000000000000001010;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule