`include "num_data.v"

module w_rom_29 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000000110001000000000010010011000000000010111011111111111011010101111111111011111100111111111101001000111111110011000010000000000101010000111111111000111001;
    mem[1] = 162'b000000001010011101111111110001010101111111110011011000000000001101110001111111111001001000000000000010000100111111111100010011111111111000011110000000000111111101;
    mem[2] = 162'b000000000000101101111111111111101001111111111111100000000000000110001010111111111100001110000000000001100011111111111111011000111111111101000000000000000001100000;
    mem[3] = 162'b111111111110110100000000000111111000111111111001001100000000000010011101000000000101100110000000000010010011111111111001000010000000000001010001111111111111110001;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111111001010111111110101010011000000000100101001111111111100110010000000000010011110000000000010011010111111111100100010000000001010101100000000000001101110;
    mem[33] = 162'b000000000000010110000000000001011000000000000001010001111111111110100000111111111110101100111111111100111111111111111011001111000000000011100010111111111011011110;
    mem[34] = 162'b111111111011011101111111111101010110111111111111001111000000000000100111000000000011001110111111111101110000111111111011110101111111111111110011000000001101101110;
    mem[35] = 162'b000000000100010000000000000011000110111111110011100011000000000100011010000000000100101101000000000010100000111111110101101101000000000000111101111111111110000001;
    mem[36] = 162'b000000000001100110000000001000010000000000000110110110000000000001110110000000000011011011111111111110100011111111111010000101111111111011011010000000000001000001;
    mem[37] = 162'b111111111100100010000000000101100100111111111001000100000000000111001010111111111001111010111111111110001010000000000000001110111111111001111001111111111011001101;
    mem[38] = 162'b000000000100111000000000000000101011111111111111100101000000000001100011000000001000010010000000001101011011000000000011101001111111111101001011000000000101110010;
    mem[39] = 162'b111111111111110011000000001000011101000000000010101000000000000101100001111111111111100001111111111011000101111111111110011111111111111110101111111111110111011111;
    mem[40] = 162'b000000000001011000000000000110000011111111111111010011111111111101111101000000000101011001111111111101111100111111111100101101000000000101101100111111110101111111;
    mem[41] = 162'b111111111101110001111111111110000001000000001000000001000000000000011100111111111010001110000000000001101001000000000110010011111111111011001100111111111110010101;
    mem[42] = 162'b000000000100011000000000000110100011000000000010011001000000000010100110111111111101001011111111111011011000000000001001111100111111110111111001000000001000001011;
    mem[43] = 162'b000000000011001100000000000110010101000000000101000011000000001000001010000000000100011111000000000010011001111111111001100110000000000010100000000000000001000001;
    mem[44] = 162'b000000000010010000111111110101010110000000000110100011000000000001110100111111111100100010000000001101010000111111110110100001000000000011110110111111111001101100;
    mem[45] = 162'b000000000010100000111111111001101110000000000001001010111111111111010011111111111111011110111111111011111110111111111110010011111111111000100100000000000000000001;
    mem[46] = 162'b000000000000110100000000000001011011111111111110100110111111110111011101111111111101010011111111111100101001000000000010111010111111111010101111000000000000001011;
    mem[47] = 162'b000000000100000011111111110111000001111111110111000101111111111111110001111111111110000101000000000001011010111111111110010011000000000000101010000000000000100010;
    mem[48] = 162'b000000000101000000000000000000000011111111111000001110111111111111000110111111111110111000111111111111000011000000000000111010111111111110101010111111111110101011;
    mem[49] = 162'b111111111100110000000000000010110010111111111110101010000000000011010110111111111000110100000000000111110110000000000100101111111111111001000011111111111110110011;
    mem[50] = 162'b000000000010011101111111111111111110111111110110000001111111110110001101000000000101001000111111111101001010111111111010010111111111111100100010000000000010101000;
    mem[51] = 162'b000000000101000100000000000110010000000000000001010101000000001010010101000000000110010000000000000011110111000000000100000011000000000001110010000000000011001000;
    mem[52] = 162'b000000000010000110000000000001101101000000000101001011000000000111111010000000000001010000000000000100111111111111111100110101111111111100110111000000000001000101;
    mem[53] = 162'b111111111110011001000000000101010000111111110001011001000000000110101011111111111101101100111111111101010111111111111101100000111111111111010111000000000011110010;
    mem[54] = 162'b111111111111110110000000000000001101000000000000101100111111111111110101111111111111110100000000000011010000000000000101010011000000000100011001000000000001010100;
    mem[55] = 162'b000000000000101000000000000010111111111111111011011100000000000010101111000000000010011100000000000001100100111111111011001110111111111011011111000000001000100100;
    mem[56] = 162'b000000000100001101111111110100001011000000000100100100111111111100001110000000000001101101111111111100110111000000001100110010111111111101000011111111111001001101;
    mem[57] = 162'b111111111101110101000000000011101001000000000110101111000000000100101110111111111001110010111111111101000010111111111111001110111111111111000100111111111001100111;
    mem[58] = 162'b111111111111010000111111111101110100000000000100011011000000000101010110000000000010011001000000001010100010000000001000111001111111110110001010000000000111001111;
    mem[59] = 162'b000000000010101001111111110111000000000000000001101010000000000010010010111111111111000111000000000011110111111111110111001101111111111110101010000000000110101011;
    mem[60] = 162'b111111111101101110000000000000001011111111111100101100000000000110110100111111111000100010000000000000111110000000000000001011000000000001010101000000000010011111;
    mem[61] = 162'b111111110110000010000000000101010011111111111111100001000000000010011100111111111001001000111111111011101001111111111100010100000000000000001101000000000001010110;
    mem[62] = 162'b000000000100001100111111111111111101111111111110111100000000000001111001000000000100110101111111111110100111111111111100010010000000000000110000000000000001111000;
    mem[63] = 162'b111111111011111110000000000000111000000000000000101011111111111100110100000000000101001010000000000101100101000000001001000110000000000011110101000000000000101010;
    mem[64] = 162'b111111111111111010000000000011000011000000000100000110000000000000111010000000000111000000111111111110011100000000000001101110111111110111100100111111111011111110;
    mem[65] = 162'b111111111110011100111111111010110010000000000001010001111111111100101110111111111111011100000000000000101011000000001000000101000000000100101010000000000001000110;
    mem[66] = 162'b111111111010011011111111111101001101111111111100000110000000000001100011111111111100110001000000000000011110000000000001100100000000000101111010000000000010011000;
    mem[67] = 162'b000000000110001101000000000001100100111111111101111000000000000011010111000000000000001101000000000000101111111111110110001000111111111011111111000000000000110110;
    mem[68] = 162'b111111111111100110000000000001000011000000000011101000000000000001001000000000000100001000111111111011110110000000000010001000111111111110011100111111111110101100;
    mem[69] = 162'b111111111100010111111111110111111010000000000110011111000000000011011011000000000110010101000000000001110100000000000000110001111111111111110101000000000000101010;
    mem[70] = 162'b111111111111110100000000000000110010000000000001000010000000000100011101000000000000100001000000000010111000111111110101110011000000000011000001111111111110110100;
    mem[71] = 162'b000000000100011110000000000011111110000000000011001101111111111100100100000000000100111010111111111100000111000000000101111101111111111110100111111111111100100001;
    mem[72] = 162'b000000000100100110000000000000001100111111111101001111111111111011100110000000000000000111000000000010101101111111110110111011000000000010011000000000000010110110;
    mem[73] = 162'b111111111000111110111111110001010001111111111110111001000000000100100111111111111010110111000000000100011101000000000000111101000000000000010100111111111011110000;
    mem[74] = 162'b000000000100011001111111111100001000111111111000000010111111111110100010111111111111100100000000000010011100111111111100110101111111111110001101111111111011001010;
    mem[75] = 162'b111111111001100001000000000001110011000000000110001011111111111101001010111111111000100011111111111111001010111111111110100011111111111101000000111111111111001100;
    mem[76] = 162'b000000000001110101000000000011000011000000000101001110111111111101100001000000001010101110000000000110101011111111111110000001000000000011010111000000000010111110;
    mem[77] = 162'b000000000010111101000000000010001001111111111110010010000000000010100100000000000000100110000000000001001110111111111010010111111111111000101111111111111111100101;
    mem[78] = 162'b000000000101001010000000001010101000000000000011111010000000000010101010000000000011110110000000000101111111111111111011110010000000001010100000111111111000110010;
    mem[79] = 162'b111111111000001101111111111100010101111111111110000110111111111011100001000000001000010101000000000000001001111111111101110001111111111010101110111111111100111101;
    mem[80] = 162'b000000000111100010111111111001100101111111111111000101000000000011001001000000000011011011111111111111000100111111111100000010000000000100111000111111111001110110;
    mem[81] = 162'b000000000101010101111111111011010001000000000010110101000000000000011010000000000010000011111111111011100101111111111001100010111111111111010011111111111110100111;
    mem[82] = 162'b000000000010101101000000000011100000000000001001011100111111111011110001111111111101010001000000000100111011000000000011100001000000000010100000111111111110010000;
    mem[83] = 162'b000000001001101010000000000011010110000000000101110111000000000001110101111111111101001001111111111001000001000000000110011011000000000010111010111111111001100101;
    mem[84] = 162'b111111111101100100111111111110101000111111111010011111000000000001010110000000000010001010000000000000110010111111111010001101000000000000100011000000000100101011;
    mem[85] = 162'b111111111101010011000000000101100101000000000101000111000000000111011011111111111111010001000000000010111111111111111101110100000000000011101001111111111110010000;
    mem[86] = 162'b000000000111001110111111111100101110000000000111000001000000000110001001000000000100111001000000000110010110000000000001000000000000000101001100000000001000100011;
    mem[87] = 162'b000000000010011110111111110110110100111111111111110110000000000011000101000000000011011011000000000010010110111111111010101010111111111111100110111111111110011110;
    mem[88] = 162'b111111111110100111000000000001100010111111111101001000000000000000100111111111111111111011000000000000010001111111111101000011000000000011011010111111111000111101;
    mem[89] = 162'b000000000011011000000000000010100100000000000000011110111111111110100110111111111011001110111111111111001111111111111100001000111111110111011011111111110101000110;
    mem[90] = 162'b111111111101111001000000000000100101000000000110100010111111111111001101000000000110011110000000000011001010000000001001101011111111110111111000000000000010101010;
    mem[91] = 162'b111111111111011001111111111010000111000000000111111001000000000000010100000000000000010000000000001000010101111111111100110111111111111100100001111111111101011000;
    mem[92] = 162'b000000000001001001111111111110100110000000000100010011000000000101001101111111111101110111111111110111110100111111111101000101000000000001010101111111111101010101;
    mem[93] = 162'b000000000111101100000000000000111000111111111111100111000000000011110111000000000001100011111111111101100110000000000001011011111111111110001011111111111101001101;
    mem[94] = 162'b111111110110001111000000000000010010000000000001100101111111111101100111111111111110001011000000000110011101000000000000010101000000000011011110111111111111110100;
    mem[95] = 162'b111111111101011011111111111010111111000000000011010101000000000111011100000000000001010000000000000000010010000000000110110111111111111101100010000000000000001101;
    mem[96] = 162'b111111111111101011111111111111111010000000000000010100000000000000000010000000000000000000000000000000000011111111111111110100111111111111111110000000000000010001;
    mem[97] = 162'b000000000000010110000000000000000000000000000000001001000000000000001000111111111111110100111111111111111001111111111111110011000000000000000011000000000000010100;
    mem[98] = 162'b000000000000001001000000000000000110111111111111111011000000000000001000000000000000011000111111111111110010111111111111110111111111111111111001111111111111110011;
    mem[99] = 162'b000000000000010101000000000000000101111111111111111100000000000000000010000000000000001010111111111111110101000000000000001001000000000000000001111111111111111000;
    mem[100] = 162'b000000000000001110111111111111111010111111111111111000000000000000001100000000000000000001000000000000001011000000000000000011000000000000001000000000000000010000;
    mem[101] = 162'b111111111111110001111111111111111011000000000000001010000000000000010010000000000000000111111111111111110010000000000000000010000000000000000100000000000000010100;
    mem[102] = 162'b000000000000001101000000000000001010000000000000001101000000000000000110000000000000000110000000000000001101000000000000000011000000000000001100000000000000000100;
    mem[103] = 162'b111111111111100010000000000000001011111111111111111001000000000000000001000000000000010001000000000000001110000000000000001100000000000000010001111111111111110110;
    mem[104] = 162'b111111111111101100000000000000000000000000000000010111111111111111110001000000000000000000111111111111111110000000000000000101000000000000001000000000000000010000;
    mem[105] = 162'b000000000000001011000000000000001011111111111111111001000000000000001100000000000000000100000000000000000010000000000000001111111111111111111110111111111111110110;
    mem[106] = 162'b111111111111111011000000000000001000000000000000001000111111111111111100000000000000000111111111111111111011111111111111111010000000000000001000111111111111111110;
    mem[107] = 162'b000000000000000100111111111111110011000000000000000110000000000000000110000000000000000100111111111111111100111111111111110011111111111111111010111111111111110000;
    mem[108] = 162'b111111111111110010111111111111111111111111111111110100000000000000000011000000000000001100000000000000010011000000000000000010111111111111111101111111111111111010;
    mem[109] = 162'b111111111111111100111111111111101001000000000000000100111111111111111100111111111111111100111111111111111011000000000000001011111111111111111101111111111111110000;
    mem[110] = 162'b111111111111110111000000000000010000111111111111110001111111111111111100111111111111111100111111111111111011000000000000001011000000000000000101000000000000001101;
    mem[111] = 162'b000000000000001101000000000000000010111111111111111010000000000000001010111111111111111111111111111111101001111111111111111000000000000000001011111111111111110111;
    mem[112] = 162'b000000000000010100000000000000000111000000000000011100000000000000000110111111111111111001000000000000000100000000000000110110111111111111101111111111111111101110;
    mem[113] = 162'b000000000000010110111111111111111011111111111111110100000000000000000001000000000000001010111111111111110010111111111111110011000000000000000100111111111111110111;
    mem[114] = 162'b000000000000011010111111111111110100000000000000010101000000000000000110000000000000000100000000000000000111000000000000000011111111111111110011111111111111100001;
    mem[115] = 162'b000000000000000011111111111111110111111111111111110101000000000000000011000000000000010010111111111111111111111111111111111011111111111111110100111111111111100101;
    mem[116] = 162'b000000000000010010000000000000000000000000000000001101111111111111111001111111111111110110000000000000100110000000000000001100000000000000000111111111111111110100;
    mem[117] = 162'b000000000000001111000000000000000000111111111111100100000000000000001010111111111111110010000000000000010000000000000000001100111111111111101011111111111111100110;
    mem[118] = 162'b000000000000001101000000000000010010111111111111110100111111111111100110111111111111111100000000000000000000111111111111111001000000000000001011000000000000010000;
    mem[119] = 162'b000000000000001111000000000000000011000000000000010000000000000000010001000000000000010001000000000000001101000000000000001010000000000000010011000000000000001001;
    mem[120] = 162'b000000000000000110111111111111101101000000000000010011000000000000000000111111111111111101000000000000001010000000000000001001000000000000000001111111111111111101;
    mem[121] = 162'b000000000000000001111111111111101111111111111111110111000000000000000101000000000000000000111111111111110101111111111111111110111111111111111110000000000000110111;
    mem[122] = 162'b000000000000010001000000000000000001111111111111110101111111111111111010000000000000001100000000000000000110000000000000001011000000000000000101111111111111110110;
    mem[123] = 162'b111111111111100010111111111111100110111111111111101010111111111111101111111111111111111101000000000000000100111111111111101101000000000000000110000000000000001101;
    mem[124] = 162'b000000000000010100000000000000010001000000000000001011111111111111111011111111111111111001111111111111111101111111111111111111000000000000000000000000000000000100;
    mem[125] = 162'b000000000000000100111111111111111110111111111111111001000000000000000011000000000000001010000000000000000101111111111111111100111111111111110110111111111111111001;
    mem[126] = 162'b111111111111110101111111111111011111111111111111101011111111111111101111000000000000010000000000000000000100111111111111110001111111111111111110111111111111111010;
    mem[127] = 162'b111111111111111111000000000000001000000000000000001001000000000000010111000000000000001001000000000000000101000000000000001000000000000000000101000000000000001001;
    mem[128] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[129] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[130] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[131] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[132] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[133] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[134] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[135] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[136] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[137] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[138] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[139] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[140] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[141] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[142] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[143] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[144] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[145] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[146] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[147] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[148] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule