`include "num_data.v"

module w_rom_10 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b111111111010010011111111111011100101000000001010001010000000000101111100000000000010101010111111111011101101111111111111110011000000000110110000111111111011000000;
    mem[1] = 162'b111111111101101011111111111111100001000000000101000110111111111100101110111111110100001101000000000111001000111111111010111010111111111110010011111111111110001011;
    mem[2] = 162'b111111111100010001111111111111101011000000000011010000111111111101011011111111111110000110111111111100000111000000000110110000111111111000110111000000000000001100;
    mem[3] = 162'b000000000111010111000000010110001110111111101001110101000000001000110101111111101111101011000000001001110011111111110110100101111111111101011110111111110100110110;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111110110110010111111111111101110111111111110111010000000000101011010111111111111100011111111110110010010000000000100011101111111111110101001000000000101001110;
    mem[33] = 162'b000000000101001000111111111101110110000000000110010100111111111111010010111111111101110100000000000100010100111111110011000000111111111111110010000000000001111100;
    mem[34] = 162'b000000000000111110111111111100100000111111111000000010000000000001111001111111110111011100111111111100000000000000000011000101000000000001110111000000000011110001;
    mem[35] = 162'b000000000001011000111111111100011010111111111111011110000000000100100011000000001010000001111111111100111110000000000101011011000000000101100000111111111100111111;
    mem[36] = 162'b111111111101110000000000000001001110111111110111010000000000000110111110111111111110100100111111111111101010000000000000001111000000000101000100111111111100100000;
    mem[37] = 162'b111111111001110111000000000000100001000000000100010100000000000011011100000000000011000011111111111000110110111111111111100000111111111001000100111111110111010010;
    mem[38] = 162'b000000000111100111000000000101101100111111111111001011111111111101001011000000000110001111000000000010101011000000000101011010000000000101001110000000001000011110;
    mem[39] = 162'b111111111110000011000000000000000011000000000010010101111111110111011101111111111100101111000000000010001101111111111101101110000000000110000001000000000010010000;
    mem[40] = 162'b111111111100000111000000000011111111000000000001110110000000000000110001000000000100010110000000000100110010000000000001110101111111111011011011000000000010111000;
    mem[41] = 162'b111111111011110101000000000100011010111111110101101001111111110111100000111111111101010111000000000000100110000000001001110011111111111011001000111111111000001111;
    mem[42] = 162'b111111111011100000000000000000000011000000000000111001111111111111000010111111111110100000000000000010111100111111111011111001111111111011111101111111111011010001;
    mem[43] = 162'b111111111110110101000000001010010111111111111110000110000000000000010100111111111111110100000000000010111011111111111001000111000000000011011010000000001000101001;
    mem[44] = 162'b000000000000100000111111111100111000000000000011010100111111111111100011111111111111111100111111111100001111000000000111011111111111111101101001111111111011111100;
    mem[45] = 162'b000000000000011000000000000010000010111111111110001101111111110111111100111111111110111010111111110110011111000000000010101111111111111010111101000000000011011010;
    mem[46] = 162'b000000001000001010000000000110001111111111111111110111111111111000100001000000000001000011111111111111100110111111111101110011000000000001110010111111111001110010;
    mem[47] = 162'b000000000100100011000000000110110001111111111100010010111111111101010001111111111101111000111111111010000010000000000100110010000000000011011100111111111011010000;
    mem[48] = 162'b000000000110110110111111110110100101111111111011110011111111111100000000000000000001001001111111111110010000000000000111000111000000000110111001000000000001001001;
    mem[49] = 162'b000000000011101001000000000000001010000000000011111100000000000010001110111111111101001111000000000000100011000000000100111000111111110101011110111111111101111110;
    mem[50] = 162'b000000001000111101111111111011100011111111111111111011111111111101001001000000000000000011111111111111001011111111110110110000000000000000110111000000000001011100;
    mem[51] = 162'b000000000001011101000000000011111000111111111101100000000000000011001010000000000100011100111111111101000101000000001000101010000000000101101011111111111111111100;
    mem[52] = 162'b000000000111100101111111111100110001111111111100110011000000000110011011000000000110001001000000000111000100111111111111101101000000000101010100000000000001101110;
    mem[53] = 162'b111111111101101101111111111101001011111111111111100010000000000000010011111111111011001000000000000010111100111111110010111011000000000011001000000000000001000101;
    mem[54] = 162'b111111111101111111111111111101000011111111111101111011111111111110010111111111111110110001000000000001000010000000000000001110000000000100000111000000000110100001;
    mem[55] = 162'b000000000110000101111111111001010011000000000111110001000000000000010000000000000001111111111111111100110111111111110001010001111111111110111000111111111100001000;
    mem[56] = 162'b000000000011010111111111111110110011000000000000000001111111111110001101000000000100010010111111110111011011000000000010001000000000000101011111111111110011101000;
    mem[57] = 162'b000000000010001000111111111101110001000000000011001001000000000100000011111111111101001111000000000000100101000000000101011000111111111001101110000000000101101101;
    mem[58] = 162'b000000000010001110111111111111111000111111111010101111111111111111100100000000000101110010111111110111011010000000000001000011111111111000110011000000000001110100;
    mem[59] = 162'b111111111110010000000000000001010011111111111100011010000000001010001001000000000101000011111111111110110000111111111001101010111111111111100101111111111101111111;
    mem[60] = 162'b000000000010111000000000000000101111000000000110001111111111111111000110000000000011010001111111111010011110111111111101001000111111111110001011111111111110110011;
    mem[61] = 162'b000000000011101100000000000011101110111111110101110101111111111101100100111111111101111011000000001001101000111111111010010000111111111101111000000000001000111010;
    mem[62] = 162'b111111111101101101111111111110001110111111111110000001000000001001011001111111111100111011000000000100111100000000000101000111000000000000011101111111111110011111;
    mem[63] = 162'b000000000100011110000000000001101101000000000100001010000000000011101011111111111101000101111111111111001010000000000010110101000000000001111110111111111101000100;
    mem[64] = 162'b000000000100011101000000000100110101000000000001010110111111111110100101000000000010110110111111111000010110000000000010101001000000001011001101111111111001100001;
    mem[65] = 162'b000000000000101100111111110111111010111111111110010100111111111111110101000000000010001001000000000101011011000000000111000010000000000000010001000000000000100111;
    mem[66] = 162'b000000000001001101111111111101011001111111111101100101111111111110011111000000000000101001111111111110110101000000000010011110000000000000111111000000000010100101;
    mem[67] = 162'b000000000010110111111111111100011100111111111111101101111111111110101100111111111010111011000000000010110111000000000001000101000000000010001110111111111100101001;
    mem[68] = 162'b000000000001011010000000000101001010000000000000100001111111111010010111111111110110000110000000000111011000111111111100101000111111111101111100000000000010101100;
    mem[69] = 162'b000000000000001100111111111111011000000000000010110100111111111100100101111111111100111101000000000000011011111111111010010000111111111111100001000000000100011101;
    mem[70] = 162'b000000000001101000000000000001101011000000000001000010000000000011000110000000000000011111000000000001000001111111111110100111111111111111110001000000000000110110;
    mem[71] = 162'b000000000111100100000000000001110000000000000100001001000000000010101011000000000110011000111111111011111010111111111011111010000000000111001111000000000001111010;
    mem[72] = 162'b000000000011001100000000000011011000000000000000110111111111111110101101111111111110000000111111110101001001000000000001111000000000000000001010111111111100110010;
    mem[73] = 162'b000000000011100101000000000000101011111111111101111001000000000000001011111111111001100111000000000100010010111111111110110011111111111010100011000000000010010100;
    mem[74] = 162'b111111111001111000111111111111110101000000000010011110111111111110000110000000000001111000111111111111101001000000000011011000111111111110101110000000000101111111;
    mem[75] = 162'b111111111110000001111111111011000010000000000001011011000000000100101100000000000000110000111111111100101000111111111011001101000000000101000110111111111111100000;
    mem[76] = 162'b000000000010110110111111111100100111111111111111101011000000000010100011111111111111110010000000000100101011000000000001101110000000000010111110111111111111010011;
    mem[77] = 162'b111111111100111101111111111100101010000000000100010101000000000000000000000000000000101010000000000101110100000000000010000101000000000100111100000000000000011110;
    mem[78] = 162'b000000000001100101000000000001010101000000000101001111000000000010010100000000000100001101111111111101110111000000000010000100000000000110011101111111111111101111;
    mem[79] = 162'b111111111100010000000000000010101000000000000100001101111111111100111100000000000010000110000000000000110110000000000001101011000000000011010000000000000101011100;
    mem[80] = 162'b000000000010100010111111111110100101000000001000000011111111111100000011000000000001000011000000000010100010000000000011010111000000000001101011000000000101010001;
    mem[81] = 162'b000000000000001001111111111111101000000000000001111100111111111111000010000000000000000001111111111100101100000000000000010001111111111111111010000000000000010010;
    mem[82] = 162'b111111111010010100111111111111110010000000000100011001000000000100111000000000000010010111111111111001101001000000000111001100000000000100101101111111111110011011;
    mem[83] = 162'b111111111110010111000000000101001100000000000001101010000000001000011000111111111101110100111111111010011000111111111100110010000000000110101011111111111101111100;
    mem[84] = 162'b000000000001100010111111111110000011000000000100010111111111111011010100111111111101100111111111111110000101111111111100011111111111111111001001000000000111011011;
    mem[85] = 162'b111111110111010011000000000010011111000000000110010111000000001000100000111111111110000111000000000001001001000000000000101101000000000000111110111111111111111001;
    mem[86] = 162'b111111111111101011000000000101011000000000000111011000000000000100110110000000000100100001000000000101101001000000000000001101000000000110001000000000000000110000;
    mem[87] = 162'b000000000011111111111111111101110101111111111010110110000000000110111010000000000011000100111111111101110110000000000111101001111111110110111110111111111101010111;
    mem[88] = 162'b000000000011010101111111111110000101111111111111010010111111111111011001111111111101110000000000000100000011000000000001000000000000000010101111000000000011000010;
    mem[89] = 162'b111111111001110111111111111011011001000000000101110011000000000001010010111111111011111100000000000011001011111111111110100110000000000111101010111111111011101110;
    mem[90] = 162'b000000000101000111000000000100110100000000000001111111000000000110110001000000000010101100000000000001010110000000000000010101000000000000000011111111111001010010;
    mem[91] = 162'b000000000001011000111111111111101010000000000110110100111111111100011010000000000010000011111111111110110110000000001001110111000000000101101010111111111011010010;
    mem[92] = 162'b000000000010000011111111111100010010111111111101100110111111111111111010111111111100111011000000000000001110111111111111010000111111111111011011000000000001101010;
    mem[93] = 162'b000000000000010000000000000001101110000000000010111100111111111100001010111111111011000001000000000100111100111111111001101110000000000001110111000000000101101101;
    mem[94] = 162'b111111111110011000111111111110100000000000000010000011111111111101110000111111111110010111000000000010101110111111111111010111000000000001001011000000000100100001;
    mem[95] = 162'b000000000000110111000000000111111000000000000100000001000000000010011010111111111101111100000000000000110011000000000001000100000000000000001100000000000001100001;
    mem[96] = 162'b000000000000000101000000000000001001111111111111111111000000000000010110111111111111111100111111111111111000111111111111100111111111111111100101000000000000000100;
    mem[97] = 162'b000000000000010101111111111111110101000000000000000101000000000000010111000000000000000011000000000000001000111111111111101001111111111111110111000000000000000001;
    mem[98] = 162'b000000000000001010111111111111111110111111111111111110000000000000001000000000000000001000111111111111111000111111111111100101000000000000001011111111111111101010;
    mem[99] = 162'b000000000000100110000000000000011110111111111111111001000000000000001100111111111111111001111111111111110010000000000000000011111111111111111101111111111111101100;
    mem[100] = 162'b111111111111110111111111111111101011111111111111111000000000000000000110111111111111110011000000000000001001111111111111111101000000000000000000000000000000001111;
    mem[101] = 162'b000000000000010110000000000000001010000000000000000000000000000000000001111111111111101011111111111111110011111111111111101011000000000000000101000000000000000000;
    mem[102] = 162'b000000000000010001000000000000001110000000000000000101111111111111101101111111111111101110111111111111101101000000000000000110000000000000000101111111111111111110;
    mem[103] = 162'b111111111111111100000000000000001110111111111111111101111111111111111000111111111111111011111111111111111111111111111111111000111111111111111010111111111111110101;
    mem[104] = 162'b111111111111111001000000000000000000111111111111100111111111111111101110111111111111111011111111111111110101000000000000010111000000000000001011000000000000000010;
    mem[105] = 162'b000000000000000100111111111111110100111111111111111111000000000000001111111111111111111101000000000000000001000000000000001100111111111111101100111111111111110011;
    mem[106] = 162'b111111111111111100000000000000000000000000000000000100111111111111110001111111111111101101111111111111111111000000000000000101111111111111110010111111111111110100;
    mem[107] = 162'b111111111111111110111111111111111011000000000000000011111111111111111111111111111111111011111111111111111000111111111111111011111111111111111001111111111111111010;
    mem[108] = 162'b111111111111111011111111111111111110111111111111101111111111111111101000111111111111101101000000000000000010111111111111101111111111111111101111000000000000000010;
    mem[109] = 162'b111111111111101000111111111111111001000000000000001100000000000000000011111111111111111110000000000000000100111111111111111000111111111111110011000000000000000000;
    mem[110] = 162'b111111111111111101000000000000001100111111111111111011111111111111111001000000000000000001111111111111111001000000000000001011000000000000000101000000000000011001;
    mem[111] = 162'b000000000000000110111111111111111101000000000000000000000000000000001101111111111111111001111111111111100111111111111111111000000000000000000011111111111111110011;
    mem[112] = 162'b111111111111111001111111111111111111000000000000011111000000000000001101111111111111110100111111111111110111000000000001011001111111111111101110000000000000001111;
    mem[113] = 162'b000000000000001111111111111111111001111111111111111111111111111111110111000000000000000110111111111111110000000000000000010010111111111111111101000000000000000100;
    mem[114] = 162'b000000000000001010111111111111110100111111111111011010000000000000000011000000000000000000000000000000001100000000000000000110111111111111111010111111111111101010;
    mem[115] = 162'b111111111111111111111111111111111101111111111111111001111111111111110010111111111111111101111111111111111110111111111111111011111111111111111000000000000000000001;
    mem[116] = 162'b000000000000000000111111111111111010000000000000010101000000000000011011000000000000000110000000000000001001000000000000010010000000000000001001111111111111111100;
    mem[117] = 162'b000000000000000100000000000000000100111111111111101100111111111111110011111111111111110111000000000000000000111111111111111010111111111111101000111111111111110001;
    mem[118] = 162'b000000000000000011111111111111111111000000000000000001111111111111100010111111111111100110111111111111110000111111111111111111111111111111111111111111111111111011;
    mem[119] = 162'b000000000000001111000000000000000110000000000000000000000000000000010110000000000000001010111111111111110110000000000000001111000000000000010010000000000000001100;
    mem[120] = 162'b111111111111110110000000000000000001000000000000001100000000000000000010000000000000001010000000000000000001111111111111110110111111111111111000111111111111111111;
    mem[121] = 162'b111111111111110010111111111111110110111111111111101000111111111111110110111111111111111000000000000000010111111111111111100100000000000000010100000000000000010001;
    mem[122] = 162'b000000000000001011000000000000000111000000000000001101000000000000000000111111111111110001000000000000000011000000000000010101111111111111110110111111111111110111;
    mem[123] = 162'b111111111111100001111111111111101101111111111111111010111111111111110100111111111111110101111111111111111110111111111111111010000000000000000011111111111111111011;
    mem[124] = 162'b000000000000010011000000000000011000000000000000000010111111111111111110111111111111110100111111111111111001000000000000001010111111111111110011111111111111111110;
    mem[125] = 162'b111111111111111111000000000000000010111111111111111100111111111111111110000000000000000110111111111111111100111111111111110100111111111111110100000000000000001100;
    mem[126] = 162'b111111111111110011111111111111110110111111111111111100111111111111111110111111111111101100000000000000001000111111111111110110111111111111111101000000000000000011;
    mem[127] = 162'b111111111111101010111111111111110110111111111111110101111111111111111100111111111111110001111111111111101100000000000000011000000000000000001010000000000000010100;
    mem[128] = 162'b111111111111111011111111111111110101111111111111101001000000000001010011111111111111100101111111111111100000111111111111000111111111111111111111111111111111011101;
    mem[129] = 162'b111111111111111101111111111111111010111111111111110011111111111111111101000000000000000001111111111111111001000000000001001010111111111111110100000000000000001000;
    mem[130] = 162'b000000000000000101111111111111111000111111111111111010111111111111110110111111111111111110111111111111111100111111111111111100111111111111111000111111111111111100;
    mem[131] = 162'b000000000000000111111111111111111101000000000000000010000000000000000000111111111111110001111111111111110000111111111111111100111111111111111101111111111111111011;
    mem[132] = 162'b000000000011011000000000000000111000000000000010010010000000000011010111000000000001011001111111111111100111111111111111111011000000000000010000000000000000001000;
    mem[133] = 162'b111111111111111011000000000000000000000000000000000111000000000000000101000000000000000000111111111111111011000000000000011100000000000011110011000000000100001110;
    mem[134] = 162'b111111111111110011000000000000000010111111111111101111000000000000001000111111111111111101000000000000000100111111111111111101000000000000000111000000000000000100;
    mem[135] = 162'b000000000000011001000000000000011011111111111111110010111111111111110100000000000011010111000000000000000000000000000000010010111111111111111011000000000001100110;
    mem[136] = 162'b000000000001110101000000000001110011111111111111101111000000000000001001000000000001100010111111111111011110111111111111110000111111111111101000000000000001011110;
    mem[137] = 162'b111111111111110110111111111111110101111111111111111000000000000000000001111111111111111000111111111111111111000000000100010100000000000100011000000000000100111001;
    mem[138] = 162'b000000000000000111111111111111000010111111111111010010111111111111110010111111111111101101111111111111110100111111111111110001111111111111110100111111111111110101;
    mem[139] = 162'b111111111111111100111111111111101010000000000000010001000000000000010011111111111111101000111111111111111110111111111111011110000000000000000010000000000001110010;
    mem[140] = 162'b111111111111111000111111111111111101000000000000000010111111111111111001000000000000000010111111111111101111000000000000000001111111111111111010111111111111110110;
    mem[141] = 162'b111111111111111110000000000000000010111111111111110010000000000000000000111111111111111001111111111111110111111111111111101111111111111111101111111111111111101101;
    mem[142] = 162'b000000000000000101111111111111111011111111111111111000111111111111111110111111111111111101000000000000000001111111111111110011000000000000000010000000000000000000;
    mem[143] = 162'b000000000000000001111111111111111101111111111111110010111111111111111010111111111111111100111111111111110111111111111111110111000000000000000000111111111111110100;
    mem[144] = 162'b111111111111110000111111111111111001000000000000000011111111111111110111111111111111111100111111111111111010000000000000000100111111111111110010000000000000000000;
    mem[145] = 162'b000000000000000101000000000000001000000000000000000100000000000000001101111111111111111100111111111111110011111111111111111010111111111111110110111111111111110000;
    mem[146] = 162'b000000000000000001111111111111111101111111111111111011000000000000000110000000000000001011000000000000000101111111111111111000000000000000000110000000000000000111;
    mem[147] = 162'b111111111111111101111111111111110111111111111111111010000000000000000000111111111111111110111111111111110100111111111111111001000000000000000010111111111111111110;
    mem[148] = 162'b111111111111111111000000000000001000000000000000000100111111111111110010111111111111111100000000000000000011111111111111111001111111111111111000111111111111111010;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111111111111111011111111111111111001;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule