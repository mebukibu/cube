`include "num_data.v"

module w_rom_4 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b111111111111101001000000000000010101000000000111001110111111111100111101111111111111100101111111111111010001111111111010010000000000000011101000111111111100000101;
    mem[1] = 162'b000000000111001001000000001101101001000000000011010000111111111110110101000000000010000110111111111100100100000000000110100111111111111110111010000000000001100110;
    mem[2] = 162'b111111111111110100000000000000100010000000000011111101111111111100101000111111111110111100111111110111110111000000000010110010111111111000100000111111111110100110;
    mem[3] = 162'b111111011001100100111111100100100001111111101000000110111111100100101110111111001001100100111111110001011010111111111011100101111111011100111001111111010101010111;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111110110010000000000001011000111111111100110000111111111000101000111111111001011000000000000101001011000000000101001100111111111100000000000000000111011110;
    mem[33] = 162'b111111111110101101111111111011010101000000000111110001111111111110010101111111111111010111111111111100101010111111110110100010111111111010111000000000000100101001;
    mem[34] = 162'b000000000011001100000000000001100111111111111100001010111111111110011010000000000011011011111111111111010101111111111110011111111111111011100110000000000011000000;
    mem[35] = 162'b111111111011010010000000000110100010111111111011001110111111111011100100000000000001101100111111111001011001000000000000000111000000000001111011111111111100110011;
    mem[36] = 162'b000000000100000010111111111101101110000000000101001000000000000000001000000000000011010001000000000011001110000000000000010101111111111001101111000000000001100010;
    mem[37] = 162'b000000000011010000000000000000011010111111111111000001000000000001110101000000000100011000111111111101011101111111111110001111111111111001011111111111111101001010;
    mem[38] = 162'b111111111101001001000000001000010110000000000001110000000000000010100110000000000100111100000000001100000100111111111110011000000000000010001101000000000011110001;
    mem[39] = 162'b000000001001000010000000000110010010111111111101011111111111111111110011111111111100001100111111111011011010111111111000100101000000000100101000000000000011011111;
    mem[40] = 162'b000000001001011100000000000001101110000000000011101101111111111101000001000000000010110000000000000010110111111111110111101000111111111100110001000000000011010001;
    mem[41] = 162'b000000000100100100111111111101011110111111111111011010000000000100101100000000000000110101111111111100101000111111111010101011111111111010000110111111111100101100;
    mem[42] = 162'b000000000001000000000000000001101100111111111101010000111111110111111100000000000010011100111111111110101010111111111110100100000000000000111010111111110110111101;
    mem[43] = 162'b111111111010001001000000001001001101000000000100110001000000001001010101000000000111000001000000000001000101000000000010011111111111101110011111000000000001101111;
    mem[44] = 162'b000000000100011110000000000000010111111111111110011110000000000011101010000000000011100011111111111110110110111111111010110011000000000010010110111111111010111000;
    mem[45] = 162'b111111111011011100111111111011010101111111111110110101000000000010011001000000000110001011111111111111101001111111111001100010000000000001110111111111111110010001;
    mem[46] = 162'b111111111100001110111111111010010111000000000011101010000000000110010000111111111001101011111111111000010101111111110111001100000000000110010101000000000001100110;
    mem[47] = 162'b000000000010000011111111111010001010111111111000011100000000000101101110111111111011111011000000000000110110111111111101011100111111111001100100000000000000101101;
    mem[48] = 162'b111111111001111000000000000001101011111111111111101100111111111010101011000000000010110110111111111100110110111111111101011000000000000001000110000000000110000100;
    mem[49] = 162'b111111111101100110111111111101111000000000000101000000000000000000110010000000000100101110111111111011110010111111111110111011111111111110111110111111111101100110;
    mem[50] = 162'b111111111101010100000000000001001010000000000010101000111111111111111010000000001000110101111111111010111010111111111101101101000000000011000111000000000000010011;
    mem[51] = 162'b000000000011100110000000000011101100111111111110000000000000000010100001000000000101000111000000000001100101000000000101100001000000001000000110000000000011011000;
    mem[52] = 162'b000000000000101110000000000001101010000000000010010011000000000101011100000000000100101110111111111111100111000000000000101000111111111101001110111111111101010111;
    mem[53] = 162'b111111111111010110000000000001100010111111111111000100111111111101001010111111111100010001000000000101100000111111111110101111111111111001100011111111111011101010;
    mem[54] = 162'b111111111110101101000000000011010101111111111000100111111111110101001100000000000000010010000000000011011110000000001000101101111111111010001010000000000000110110;
    mem[55] = 162'b000000000001110101000000000011011000000000000010011001000000000101101101000000000101100001000000000010000001000000000010011100111111111011100101111111111100110111;
    mem[56] = 162'b111111111101110000000000000011001101000000000011100001111111111111010000000000000110010110111111111010100100111111111101101101111111111010000011000000001000101001;
    mem[57] = 162'b111111111011111100000000000000011100000000000111010000111111111110000000000000000010001000111111111111001000000000001000100111111111111100100001000000000001000101;
    mem[58] = 162'b000000000011101000111111111111111110111111111011001101000000000101100001000000000011101101000000000011010010111111111100111010000000000011100010111111111100100000;
    mem[59] = 162'b111111110101111110000000000100111110111111111101000000000000000101000010111111110101000001000000001010010001000000000011010001111111111110011100111111111010010001;
    mem[60] = 162'b000000000100101110000000000011010010111111110010101100111111111100101101000000000110000000111111111110101100111111111011110000111111111111001101111111111110111101;
    mem[61] = 162'b111111111100101111111111111110001111000000000000101110000000000111001001111111111110101000000000000000011000111111111100110011000000000110111011111111111010100111;
    mem[62] = 162'b000000000011111100111111111110001011000000001010011000000000001101100111000000000000001011111111111100101110111111111111101011000000000010001111111111110001110011;
    mem[63] = 162'b000000000000001011000000000110110100000000000001110011000000000010100100111111111101110111111111111101101011000000000011010101000000000100111111000000000010101100;
    mem[64] = 162'b111111111011001010111111111000100111111111111011011110000000000000000001000000000001111101000000000011001110111111111110000100000000000010110000000000000001001010;
    mem[65] = 162'b111111111011000000111111111100000011111111111110110100000000000010001110111111111110100110000000000011100001000000000011110111000000000001011110000000000000111011;
    mem[66] = 162'b000000000000101010111111111100101010111111111001011000111111111011111101000000000000111010111111111011011111111111111111001011000000000011010000111111111110010010;
    mem[67] = 162'b111111111001100000111111111011011000111111111110001011000000000010101010000000000011101110000000000011110001000000000100100110111111111100100110000000000010000101;
    mem[68] = 162'b000000000001011001111111111101000110111111111101001010111111111100001010111111111010110100111111111001100110111111111100001011111111111110110000111111111010010001;
    mem[69] = 162'b111111111101011010111111111110110000000000000001101101111111111011011111111111111101000110000000000001010101111111111101011100111111111101100110111111111111110001;
    mem[70] = 162'b000000000001100001111111111111101100111111111101000010111111111011110101000000000100001101000000000011111111000000000010010000111111111101010101111111111011101010;
    mem[71] = 162'b111111111111000111111111111110111100000000000100001000000000000000111101000000000001001001111111111111000001000000001000010000000000000011010100111111111110100011;
    mem[72] = 162'b000000000011011101111111111111001101111111110111110011111111111011101011111111111110011111111111111011001110000000000001110101111111111110011101111111110111111110;
    mem[73] = 162'b111111111101111001111111111001100000111111110110000000111111111100110101111111111010011000111111111001101010111111111111111010111111111111111110111111111100001111;
    mem[74] = 162'b000000000101111010000000000001001001111111111001101010000000000010111001111111110111010001111111111110000100111111111101110000000000000001010011000000000010100011;
    mem[75] = 162'b000000000101000001111111111101110101000000000001001100000000000001110101000000000000111010000000000010011100111111111011001110000000000011101000000000000000111111;
    mem[76] = 162'b000000000001100111000000000101001101000000000010011110000000001001000011000000001101010111000000000110011010000000001100011100000000001010100111000000001001101110;
    mem[77] = 162'b000000000001000111111111111100000001000000000001001110111111111010001111111111111000111111111111111010110011111111111001100010111111111101101110111111111101100110;
    mem[78] = 162'b000000000101111011000000000111011101000000000101010011000000001001101111000000001110010111000000000101111110000000001000101100000000001000001010000000001001010011;
    mem[79] = 162'b000000000000001011111111111110011101000000000101011101000000000011100101111111111110111101000000000000001010000000000001110111111111111111111001111111111100100111;
    mem[80] = 162'b000000000011111000111111111010110010111111111000010001111111111110001011000000000000001010111111111101111000111111111101101111111111111111111011000000000000001011;
    mem[81] = 162'b000000000110011100111111111111101010111111111111001111111111111000101100111111111111001010111111111011101010111111111011001101111111111011010011000000000100101011;
    mem[82] = 162'b111111111110101000000000000100001011000000000001100010111111111101010111000000000010110100111111111010010010111111111000010101111111111011101011000000000001011100;
    mem[83] = 162'b111111111111101010111111111111110101111111111110010101000000000010011101111111111101111000000000000010111010111111111011101110000000000100011101111111111101111101;
    mem[84] = 162'b111111111111110001111111111110111111111111111001001110111111111110011110111111111111010110111111111110100111000000000100101111111111111110011001000000000101100111;
    mem[85] = 162'b111111111011110111111111111101001101111111111101100011000000000010111000000000000011100111000000000010111111000000000100011001000000000010110101000000000011101000;
    mem[86] = 162'b000000000101100000000000000010110101000000000010100110000000001001001011000000001000110100000000001001001011000000001010001110000000001101010100000000001110110110;
    mem[87] = 162'b000000000000101111111111111100101001111111111000011000000000000010110011000000000011100011111111111101011111000000000000100010111111111110101110000000000001010010;
    mem[88] = 162'b000000000010011010111111111110000001111111111110100100000000000000101011111111111110100000111111111101111101111111111001011000000000000010100110111111111111101010;
    mem[89] = 162'b111111111111010011111111111010111011111111111111111100000000000101001010111111111101101110111111111100001100111111110101101101000000000011010000111111111101001010;
    mem[90] = 162'b111111111111011111000000000001010100000000000011011101000000000001100110000000000011100111111111111101111001000000000000011100000000000101101101111111111101100110;
    mem[91] = 162'b000000000101100011111111111110111100000000000100000100000000000011101101000000000101010011000000000100110000000000000101110000000000000110000010000000000111010010;
    mem[92] = 162'b000000000011010011111111111001110110111111111100110111111111111111000101111111111111010001000000000001111010111111111001001001111111111110101100000000000011000100;
    mem[93] = 162'b111111111001111100111111111111001110000000000010000010000000000001110001000000000001000011000000000100101011000000000010001110111111111110110000000000000000010010;
    mem[94] = 162'b111111111010101100000000000000101111111111111010001100111111111111000100111111111101111111111111111101000111111111111110001001111111111110101100000000000011100011;
    mem[95] = 162'b111111111101010100111111111111011111000000000001101100000000000000001010111111111111011100111111111110101111000000000100110000000000000011101000111111111110000011;
    mem[96] = 162'b111111111111110100000000000000000110000000000000000100000000000000001100111111111111111011000000000000000100111111111111101110000000000000000001000000000000001001;
    mem[97] = 162'b000000000000000111111111111111101111111111111111110001000000000000010011000000000000001001000000000000000100111111111111110011000000000000000100000000000000000100;
    mem[98] = 162'b111111111111111010000000000000000110000000000000001001000000000000001100000000000000000101000000000000011111111111111111110111111111111111111000000000000000000001;
    mem[99] = 162'b000000000000001100000000000000010011000000000000000011111111111111110101111111111111110110111111111111101111111111111111100110111111111111110111111111111111111101;
    mem[100] = 162'b000000000000010010000000000000001000000000000000001000000000000000001110000000000000001010000000000000010100000000000000001011000000000000001101111111111111111111;
    mem[101] = 162'b000000000000000011111111111111111011000000000000010111111111111111111110111111111111111010000000000000000000111111111111111110000000000000001100000000000000001100;
    mem[102] = 162'b111111111111111010111111111111111100111111111111111000000000000000000111111111111111111110000000000000000000000000000000000001000000000000000011111111111111111010;
    mem[103] = 162'b111111111111110110000000000000010110000000000000001110111111111111111001000000000000001100000000000000010010111111111111101100000000000000000111111111111111101100;
    mem[104] = 162'b000000000000010100000000000000010000000000000000010000000000000000001100000000000000001101111111111111111100000000000000000111111111111111110110111111111111111111;
    mem[105] = 162'b000000000000001011111111111111111101000000000000000110000000000000001011000000000000000010111111111111101010000000000000001011111111111111110110111111111111110101;
    mem[106] = 162'b000000000000001001111111111111111101000000000000001111000000000000000111000000000000010100000000000000001000111111111111110000111111111111111100111111111111111011;
    mem[107] = 162'b111111111111111001111111111111110111111111111111111101111111111111110110111111111111111001000000000000000001000000000000010011000000000000010001000000000000010010;
    mem[108] = 162'b000000000000000011000000000000000100111111111111111110000000000000000001000000000000000101111111111111101010000000000000100000111111111111110110000000000000001011;
    mem[109] = 162'b000000000000011111000000000000000011000000000000011100000000000000000010000000000000000100111111111111111110000000000000000001000000000000001011111111111111111000;
    mem[110] = 162'b111111111111101010000000000000001011000000000000001111000000000000010001000000000000010011000000000000010001111111111111110001000000000000010001000000000000010010;
    mem[111] = 162'b111111111111111000111111111111111010000000000000010111111111111111111111000000000000000101000000000000010011111111111111110111000000000000001101000000000000000101;
    mem[112] = 162'b000000000000011110000000000000011001000000000000011110000000000000100011000000000000001101000000000000100110111111111111111011111111111111111111000000000000100100;
    mem[113] = 162'b111111111111111100000000000000000111000000000000000111111111111111111111000000000000000110000000000000000110111111111111110001000000000000001000000000000000110000;
    mem[114] = 162'b000000000000010011000000000000010000000000000000000010111111111111111110000000000000001101000000000000001010000000000000000100000000000000000011111111111111111111;
    mem[115] = 162'b111111111111110101111111111111111000000000000000001101111111111111110010000000000000001101000000000000001010000000000000010010000000000000001101000000000000000011;
    mem[116] = 162'b000000000000000011111111111111111100000000000000000001111111111111110000111111111111111001000000000000000011111111111111101000000000000000000010000000000000001011;
    mem[117] = 162'b000000000000000000111111111111111011111111111111100001000000000000001011111111111111111110111111111111111011000000000000001010000000000000010001000000000000000001;
    mem[118] = 162'b111111111111101001111111111111111110111111111111111110000000000000011110111111111111101110000000000000011101000000000000001000000000000000001111000000000000000000;
    mem[119] = 162'b000000000000001011111111111111111000000000000000011101111111111111111001000000000000000010111111111111111010111111111111111011111111111111111000000000000000001010;
    mem[120] = 162'b111111111111111010000000000000000000000000000000000001000000000000001011111111111111111101000000000000001100000000000000011010000000000000001110000000000000010010;
    mem[121] = 162'b000000000000001111111111111111111001000000000000001101000000000000010100000000000000001100000000000000000101000000000000110111000000000000010110000000000000001001;
    mem[122] = 162'b111111111111111101000000000000000100111111111111110000000000000000000001000000000000000111111111111111110110111111111111111111000000000000010010000000000000001111;
    mem[123] = 162'b111111111111111111111111111111111100000000000000000100111111111111111000111111111111111000111111111111101101111111111111110100111111111111111101111111111111011111;
    mem[124] = 162'b000000000000001101000000000000000001111111111111111101111111111111111111000000000000001011111111111111110010000000000000001011111111111111111001000000000000000111;
    mem[125] = 162'b111111111111110010000000000000001010000000000000000011111111111111101011000000000000000010111111111111111010000000000000010110000000000000001011000000000000000100;
    mem[126] = 162'b000000000000010001000000000000001010111111111111111110000000000000100110000000000000000000000000000000001000000000000000011010000000000000010111000000000000000101;
    mem[127] = 162'b000000000000001010000000000000000110000000000000001010000000000000000100000000000000000111111111111111100000111111111111111000111111111111100101000000000000001111;
    mem[128] = 162'b111111111111000101000000000000100001000000000000011000111111111111101111000000000001011001111111111111011011000000000000100110000000000000001101111111111111000011;
    mem[129] = 162'b111111111111111100111111111111111101000000000000000110111111111111111001111111111111111011000000000000000101111111111110000101111111111111110100000000000010001000;
    mem[130] = 162'b000000000000000000111111111111111010111111111111111100111111111111111110000000000000000010000000000000000111111111111111111001000000000000000001000000000000000100;
    mem[131] = 162'b111111111111111101111111111111111100000000000000000100111111111111111010000000000000000011111111111111111101111111111111111111111111111111111001111111111111111110;
    mem[132] = 162'b000000000011101011000000000000101111000000000010100000000000000101101110000000000100001101000000000000101000000000000000011010111111111111110100000000000001000100;
    mem[133] = 162'b111111111111111000111111111111101110000000000000000101111111111111111110111111111111101101111111111111101001000000000000011111000000000101010100000000000011101111;
    mem[134] = 162'b000000000001010110111111111111100110111111111111100010111111111111100110111111111111111110000000000000000011000000000000000010111111111111111010111111111111110010;
    mem[135] = 162'b111111111111100100000000000000010000111111111111111001111111111111110110000000000010010010111111111111111101111111111111111010111111111111011100111111111111101100;
    mem[136] = 162'b000000000000111011000000000001011001000000000010000111000000000000001001000000000000101011111111111111110101111111111111111011000000000000001010000000000000001101;
    mem[137] = 162'b111111111111100011111111111111110000000000000000000000000000000000000000111111111111110000111111111111110100000000000100000101000000000010101010000000000100010001;
    mem[138] = 162'b000000000000000100000000000001000011111111111111000000111111111111101111111111111111101001111111111111101010111111111111110111111111111111110110111111111111110110;
    mem[139] = 162'b111111111110001010111111111111100011000000000001100010000000000000000100000000000000000001111111111111011110111111111111111110000000000000100100000000000010001101;
    mem[140] = 162'b111111111111111100000000000000010000000000000000001010000000000000001101000000000000001000000000000000000000111111111111111111111111111111111111000000000000000010;
    mem[141] = 162'b000000000000000100000000000000000100111111111111111010000000000000001101111111111111111101000000000000001101111111111111111000111111111111110111111111111111110111;
    mem[142] = 162'b000000000000001100000000000000000000111111111111111110111111111111111000111111111111111101111111111111111011000000000000001010000000000000000001000000000000001101;
    mem[143] = 162'b000000000000001001111111111111111100111111111111110111111111111111110110000000000000000101000000000000000100111111111111111010111111111111110011111111111111111000;
    mem[144] = 162'b111111111111111110000000000000001000000000000000000110111111111111111011111111111111111101000000000000000011111111111111111000000000000000000001111111111111110111;
    mem[145] = 162'b111111111111110011111111111111110001111111111111101110111111111111111100111111111111110111111111111111101111111111111111110011000000000000000011111111111111110011;
    mem[146] = 162'b111111111111111010111111111111110111111111111111110010000000000000000110111111111111111101000000000000000001000000000000001001111111111111111110111111111111110011;
    mem[147] = 162'b111111111111111011111111111111101010111111111111101000111111111111111100111111111111110111111111111111110000111111111111101110111111111111110100111111111111110011;
    mem[148] = 162'b111111111111111111111111111111110101111111111111110111111111111111111100111111111111110010111111111111111100000000000000000110111111111111111011111111111111110110;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111101110000000000000000100111111111111111010;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule