`include "num_data.v"

module w_rom_20 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000001001101111111110110001110000000000011001001111111111100100001000000000000011101111111111001000100111111111100100011111111111100011111000000000000000010;
    mem[1] = 162'b000000001010100010000000001101111000000000000100111111111111111101010001000000000101110000000000000010011100111111111101101101000000001000100101111111111111001010;
    mem[2] = 162'b000000000010010111111111111110110011111111111110000001000000000011010101111111101101101101111111111101110000111111111011001011111111111101001000111111110111111110;
    mem[3] = 162'b111111011011110001000000001001001001111111111011101010000000000101011110000000000000010100111111111110000101111111101100101110111111111000111101000000000101111001;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b000000000000010001000000000010011110111111111100101000000000000010011000000000000110010001111111111100111111111111111100101101000000000001001011000000000010100001;
    mem[33] = 162'b000000000001110110111111111100000101000000001000000100111111110110101100111111111101001011111111111101101000111111111010111010111111111111011111111111110100011001;
    mem[34] = 162'b111111110110001111000000000011111111000000000000100001000000000100011110000000000011000010111111110101000101111111111100000001000000000101010110000000000011000001;
    mem[35] = 162'b000000000001000011111111111111010110111111111110010100000000000010001010111111111111000010000000000101011010111111111001101011000000000011011011111111111100101100;
    mem[36] = 162'b000000000001000111111111111101010010111111111101101010000000000011100011000000000000101101111111111001011011111111111110111100000000000011010000111111111011110001;
    mem[37] = 162'b111111111110001011000000000011110100111111111100010101000000000010100111111111111101001111111111110110011110111111111010000010111111111111011101111111111111001010;
    mem[38] = 162'b000000000011001010000000000010001011000000000101101100000000001001011111000000000011010000000000000011000111000000000000011001000000000001011111000000000010100111;
    mem[39] = 162'b111111111111011101000000000110110111111111111101111101111111111111111101111111111010101111111111111100111111111111111101111101000000000001101110000000000001001011;
    mem[40] = 162'b000000000110011100000000000111000010000000000011100110000000000000110000000000000000110010000000000000000010111111111101001101000000000110001111111111110111110111;
    mem[41] = 162'b111111111101101100111111111000011000000000000001011110000000000001011000000000000101010101111111111011110010111111111110000011000000000101001100000000000101101101;
    mem[42] = 162'b000000000000000000111111111001000001000000000111010100000000000010111010111111110110111010111111111001011001000000000100101011000000000101001110111111110100010101;
    mem[43] = 162'b000000000011110100000000000010000011000000000000000001000000001000001101000000001000101000111111111110000110111111110110110010111111111000010010000000000000010011;
    mem[44] = 162'b000000000000100010111111111101011111111111111111000110111111111111000111000000000011101010111111111111101000000000000110011100111111111110111111000000001010100011;
    mem[45] = 162'b000000000101110100111111111111001001000000000010100101111111111100010001111111111001000001111111111111011101000000000000011101111111111001111011111111111011111010;
    mem[46] = 162'b111111111100000000111111111010001000111111111111001100000000000001100101111111111101001100111111111101000110000000000000101010111111111111101111111111110101110111;
    mem[47] = 162'b000000000000001000000000000010101011111111111011011010111111111111010100111111111010110011000000000000101100000000000000011110111111111110001101000000000100110010;
    mem[48] = 162'b111111111111011011111111111011001000111111111101010000111111111100110010000000000000011100000000000000001110000000000110110110000000000100110101111111111100001001;
    mem[49] = 162'b000000000010001011000000000001010101111111111111100001111111110101101010111111110101100111111111111010001111111111111110100011111111111100010001000000000111110010;
    mem[50] = 162'b000000000101101101111111111101001000000000000011001100111111110111000100111111111100110010000000000101111000111111110110011010111111111110100110000000000010011111;
    mem[51] = 162'b000000000110111000000000000101000011000000000111010000000000000001101101000000000000001010000000000101110010000000000100000011111111111110011001000000000001001000;
    mem[52] = 162'b000000000110010011000000000001101000000000000000101011000000000011111001000000000101110001000000000010001101111111111000101100111111111010001001111111111011010000;
    mem[53] = 162'b000000000000100001111111111100110110000000000010111011111111111111110010111111111101100100111111111101100101111111111100011000111111111101001110000000000010101000;
    mem[54] = 162'b111111111010001110111111111101111100000000000011011000000000000001001010111111111010000101000000000001001010111111111011111010000000000100100000000000001001000101;
    mem[55] = 162'b111111111011001010111111111100000011000000000010111100111111111110101111000000000100101010000000000010010011111111111110010011111111111110011010000000000100000000;
    mem[56] = 162'b111111111111101111111111111001011010111111111010010101000000000100110110000000000000100101111111111101001010000000000110100001111111111111011000111111111100110100;
    mem[57] = 162'b111111111000100010000000000001110010111111111110101011000000000000101110111111111101111110111111111010101010111111111100111111000000000101011011111111111011001010;
    mem[58] = 162'b111111111100011011000000000000101110000000000000001010000000000001000100000000000100100111000000001001000011000000000001011000111111111011000011000000000000000000;
    mem[59] = 162'b000000000101100100111111111100000011111111111011011001111111111101011010000000000011001110000000000011000101000000000011010100000000000001100010000000000001101001;
    mem[60] = 162'b000000000000011010000000000000001100000000000101010010000000000111011000111111110110111100111111111111010000000000000011101111111111111101111011000000000010111000;
    mem[61] = 162'b000000000010010100000000000010001001111111111001111011111111111010110010000000000010101001000000000000111001111111111110110010111111111110001011111111111110110111;
    mem[62] = 162'b000000000001001001000000000111011111111111111001100010000000001001011101000000000100111111000000001100011101111111111110000010111111111111011101000000001101011110;
    mem[63] = 162'b111111111110011111000000001000000011000000000101101011111111111111101100000000000100001000000000000011100000000000000010100100000000000010101101000000000100010101;
    mem[64] = 162'b000000000011101110111111111110000001111111111110010001111111111101110011000000000010110001111111111011100011111111111011100011111111111001001001111111110110010000;
    mem[65] = 162'b000000000000101001111111111011111111000000000000011001000000000110011110111111111101010100111111111110101000111111111101001100000000000010100010000000000011100101;
    mem[66] = 162'b000000000000111111000000000101011001111111111010000011000000000001000001111111111111111000000000000001011010000000000000001100111111111110101000000000000000111101;
    mem[67] = 162'b111111111101100011000000000100000110000000000001101010000000000010001011000000000100111101111111111100001011111111111111110101111111111010111110111111111101001101;
    mem[68] = 162'b000000000000111001000000000000001111000000000011101100000000000001110010111111111110010110111111111011111110111111111110011110000000000100010000111111111100001100;
    mem[69] = 162'b111111111111000010111111111101001101111111111100001110000000000000101010000000000001001001111111110101100111111111111111100111111111111111011010111111111101111011;
    mem[70] = 162'b000000000100001100000000000010010101000000000010101011000000000010100101111111111111000001000000000101001010111111111101100001111111111100100101000000000000001001;
    mem[71] = 162'b111111111011011011111111111110100111111111111101100100111111111101000111111111111111011100000000000001100111000000000011011010000000000000001011111111111101110110;
    mem[72] = 162'b111111111011110011000000000110010011000000000010000000111111111101101100111111111011000101111111111010110011111111111110110110111111111010000000111111111110101101;
    mem[73] = 162'b111111111111010101000000000001110100000000000011010011000000000000001101111111111111110111111111111011011010000000000111011011111111111101000100000000000011010100;
    mem[74] = 162'b000000000011101001000000000000001101000000000001100110111111111111101011000000000100111110000000000100010010111111111101011011111111111111101100111111111110001101;
    mem[75] = 162'b000000000101000111000000000000111010000000000001010001000000000001010011000000000001101000000000000101001111111111110111001101111111111100111010111111111011101101;
    mem[76] = 162'b000000000010100011000000000100010100111111111101110010000000000111010001000000000100111110000000000010110000000000000100110010000000000000011010000000000100111111;
    mem[77] = 162'b000000000011011101111111111011011100111111111010100001000000000011100011111111111110011010111111111101110111000000000001110101111111111010110000111111111110110000;
    mem[78] = 162'b000000000011111000000000000101000111000000000100010111000000000111101110000000000100001111000000000011110100000000000111000110000000000101000100111111111111110110;
    mem[79] = 162'b111111111110011111000000000010101110111111110111011000111111111101101110111111111111000000000000000000000010000000000010100011111111111100110000111111111100001000;
    mem[80] = 162'b000000000100001110111111111100101001111111111010110001000000000100110110000000000000101110111111111001111010000000000100100001111111111111000011000000000011000000;
    mem[81] = 162'b111111110101101111111111111111101101111111111011110101000000000011100101000000000000110001111111111100100101111111111101001000111111111011010110111111111111001000;
    mem[82] = 162'b000000000010001110111111111011011000000000000011000101111111111111110001000000000001001111000000000000000111000000000000110000000000000001000011111111111000100101;
    mem[83] = 162'b000000000000000111000000000011110110111111111111010110111111111111011001111111111111010111000000000101101000000000000011011110000000000010110100111111111100100110;
    mem[84] = 162'b000000000000110100000000000000101010111111111100101110000000000000010000111111111111100110111111111100001000111111110110011000111111111111000001111111111100110000;
    mem[85] = 162'b111111111111011001000000000001100000111111111101101010111111111111111011000000000100101110000000000010010011000000000100110110111111111101100011111111111111101100;
    mem[86] = 162'b000000000111111010000000000011110001000000000010001101000000000011101110000000000011010101000000000110011110000000000101110111000000000100101001000000000100110110;
    mem[87] = 162'b111111111110000010000000000001111101111111111100100110000000000000111010111111111111111010111111111101000111000000000001001010000000000010100000111111111001101011;
    mem[88] = 162'b111111111110110110000000000000110110111111111101100111111111111111011011111111110110100000111111111111000110111111111010000110111111111100001110000000000010110110;
    mem[89] = 162'b111111111110011001111111111111100101111111111000101011000000000000110011000000000001110111000000000011010001111111111011000111111111111100011010111111111100111011;
    mem[90] = 162'b000000000100011010111111111111111101000000000110000010111111111110000111000000000000111010000000000010001011000000000001011010000000000000111010000000000010000111;
    mem[91] = 162'b000000000001100101000000000101000111000000000001011010111111111101010011111111111111101010000000000011011010000000000000100111000000000100010101111111111101110011;
    mem[92] = 162'b111111111111000011000000000000101010000000000000011001111111110111110100000000000011000001111111111011111001111111111011001010000000000010110100111111111111100001;
    mem[93] = 162'b111111111011110000111111111111001101111111111101100011000000000010011100111111111110101000111111111111110111111111111111100010111111111110111101111111111111000111;
    mem[94] = 162'b111111111010101101111111111011101101000000000010100101111111111110010110111111111101101110111111111111001000111111111100001101000000000011001101111111111111010101;
    mem[95] = 162'b000000000000111111000000000010101100111111111011111111111111111110000001111111111110001100000000000011000001000000000101010111111111111011110110111111111111011000;
    mem[96] = 162'b111111111111111101111111111111110111000000000000010101000000000000001001000000000000000110000000000000010011000000000000000001111111111111101101000000000000000111;
    mem[97] = 162'b000000000000010011000000000000000110000000000000000111000000000000010001111111111111111010000000000000000011111111111111110000000000000000000111000000000000011100;
    mem[98] = 162'b111111111111110101000000000000001111111111111111101001000000000000011101000000000000011110000000000000000001111111111111110011000000000000000111111111111111111011;
    mem[99] = 162'b000000000000011101000000000000010010000000000000001011111111111111101111000000000000000101000000000000000101111111111111110000111111111111101000111111111111100111;
    mem[100] = 162'b000000000000001110000000000000010000111111111111110110111111111111111110000000000000000001111111111111111001111111111111110001111111111111101111000000000000000110;
    mem[101] = 162'b000000000000001101000000000000001101000000000000011110000000000000010011000000000000000100111111111111111100111111111111110111000000000000001001000000000000100000;
    mem[102] = 162'b000000000000001000111111111111111001111111111111110100111111111111111000111111111111111110111111111111111101000000000000001000000000000000001011111111111111111100;
    mem[103] = 162'b111111111111111101000000000000000110111111111111111000000000000000000110000000000000000000111111111111110011111111111111101011000000000000010000000000000000001000;
    mem[104] = 162'b111111111111111111111111111111111011000000000000001100000000000000010000000000000000001000000000000000010010000000000000001001111111111111101010000000000000010101;
    mem[105] = 162'b111111111111111001000000000000000011000000000000010111000000000000000100000000000000000011111111111111110110000000000000100010111111111111110111111111111111110010;
    mem[106] = 162'b000000000000001100000000000000000101000000000000010011111111111111111101000000000000000000000000000000000101111111111111101101111111111111111100000000000000001100;
    mem[107] = 162'b111111111111101010111111111111101100111111111111101101000000000000000110000000000000000001000000000000000000000000000000001011000000000000001000000000000000000111;
    mem[108] = 162'b111111111111110001000000000000001011111111111111101101111111111111111010000000000000001111000000000000000101111111111111110010000000000000000110111111111111101111;
    mem[109] = 162'b000000000000000111000000000000000001000000000000001100000000000000000000000000000000010010000000000000001000000000000000010000000000000000000101000000000000000111;
    mem[110] = 162'b111111111111111101000000000000001000000000000000000110000000000000000100000000000000000010000000000000001000000000000000000110000000000000010111000000000000000111;
    mem[111] = 162'b111111111111111111000000000000000111000000000000011101111111111111111010000000000000001001111111111111111100111111111111111000000000000000010011111111111111111100;
    mem[112] = 162'b000000000000010001000000000000001000000000000000101101000000000000010001111111111111101111111111111111110011111111111111010000000000000000011111000000000000000101;
    mem[113] = 162'b000000000000001110111111111111101101111111111111110001000000000000001110111111111111111110111111111111110100111111111111111011111111111111111111000000000000001111;
    mem[114] = 162'b111111111111111001111111111111110110000000000000001111111111111111111011000000000000000001000000000000000101000000000000001110000000000000000110000000000000000000;
    mem[115] = 162'b111111111111110100000000000000000011111111111111111011000000000000000001000000000000001000000000000000001011000000000000001010000000000000001010111111111111111100;
    mem[116] = 162'b111111111111101101111111111111110111000000000000001110111111111111100011000000000000000110000000000000000010000000000000001110000000000000000000111111111111101111;
    mem[117] = 162'b000000000000000111000000000000000001111111111111101000111111111111111111111111111111110011000000000000000111111111111111111110000000000000010001111111111111111000;
    mem[118] = 162'b000000000000010001000000000000010010000000000000000010111111111111111100111111111111101001000000000000000110111111111111111101000000000000000100000000000000010110;
    mem[119] = 162'b111111111111101011000000000000000011000000000000001100000000000000010100000000000000000110111111111111111110111111111111111000111111111111111010000000000000001100;
    mem[120] = 162'b000000000000010101000000000000000100000000000000000001000000000000000111000000000000000100000000000000011011111111111111110111111111111111101010111111111111111011;
    mem[121] = 162'b000000000000001110000000000000001111000000000000001011000000000000011010000000000000000000000000000000010000000000000001011000111111111111101001000000000000101110;
    mem[122] = 162'b000000000000001011000000000000000001000000000000000001000000000000000100000000000000000101000000000000001011111111111111111001111111111111110111111111111111110110;
    mem[123] = 162'b111111111111110111111111111111110010000000000000001011000000000000001100000000000000000000111111111111110011111111111111110110111111111111101110111111111111101101;
    mem[124] = 162'b000000000000001000000000000000011001000000000000011000111111111111110111111111111111111010000000000000000100111111111111111110000000000000010001000000000000001010;
    mem[125] = 162'b111111111111110101111111111111110000111111111111101110111111111111111111000000000000001011111111111111111111111111111111111000000000000000001100000000000000000100;
    mem[126] = 162'b000000000000010100111111111111101001000000000000010011111111111111111001000000000000000001000000000000100001111111111111110110000000000000010100000000000000001110;
    mem[127] = 162'b111111111111100010111111111111111110111111111111111010111111111111111111111111111111111101111111111111011100000000000000000100000000000000001010000000000000000101;
    mem[128] = 162'b111111111111110010000000000001111111000000000011110101000000000101100110000000000000010110111111111111010010000000000001011000000000000000000001000000000000110001;
    mem[129] = 162'b111111111111111111111111111111111000111111111111111001111111111111101100111111111111110011111111111111111110000000000000110001111111111111011010111111111111011100;
    mem[130] = 162'b000000000000000110111111111111111010111111111111111011000000000000000011111111111111110110111111111111111111111111111111111111000000000000000001111111111111111101;
    mem[131] = 162'b111111111111110100000000000000000011000000000000001000111111111111111100111111111111111110111111111111111011111111111111111000111111111111110001000000000000001101;
    mem[132] = 162'b111111111111101110000000000001000001111111111111111010111111111111111010111111111111101111111111111110111000000000000000011010000000000000111011000000000000000011;
    mem[133] = 162'b111111111111111110111111111111101101111111111111111110000000000000001011111111111111111000111111111111110110000000000000110011000000000000101101111111111111100011;
    mem[134] = 162'b000000000110001001000000000010110000000000000101010001000000000000000011000000000000000001111111111111111111111111111111111101000000000000000100111111111111110111;
    mem[135] = 162'b111111111111010000000000000000111110111111111111111010111111111111001111000000000000110010000000000010110010000000000001111000111111111111111011000000000100001100;
    mem[136] = 162'b000000000000000011111111111111111101111111111111110101111111111111111111111111111111110101111111111111111101000000000000000111111111111111111101000000000000000001;
    mem[137] = 162'b111111111111111101111111111111111100000000000000010001000000000000001010111111111111111100111111111111110110000000000000001001000000000000000110111111111111111010;
    mem[138] = 162'b111111111111111011111111111111111101000000000000000101000000000000000000000000000000000010000000000000000111111111111111110100111111111111111011111111111111101100;
    mem[139] = 162'b000000000000001100000000000000000111111111111111111101111111111111111111000000000000000000000000000000001010111111111111101111111111111111110111111111111111111110;
    mem[140] = 162'b000000000100101000000000000001010101000000000100101010000000000001110100111111111111111001000000000001000110111111111111011110111111111111110010111111111101011010;
    mem[141] = 162'b000000000000000111111111111111111100000000000000001001111111111111111110000000000000000100000000000000000111000000000011011011000000000011110010111111111111110111;
    mem[142] = 162'b000000000011010110000000000100001011000000000011101000111111111111111000111111111111111000000000000000001000111111111111111110000000000000000101111111111111111111;
    mem[143] = 162'b000000000000000010000000000000110110111111111111000111000000000001101110111111111111100011111111111111000111000000000000111011000000000001000110000000000011110000;
    mem[144] = 162'b000000000000001010000000000000000100111111111111111011111111111111111110000000000000000011000000000000010000000000000000000101000000000000001010000000000000001011;
    mem[145] = 162'b000000000000000110000000000000000110111111111111111010111111111111111100111111111111111100111111111111111001000000000000000011111111111111110101000000000000000001;
    mem[146] = 162'b000000000000010100000000000000000110111111111111110110111111111111111001000000000000000111111111111111111101000000000000000010111111111111111001111111111111111001;
    mem[147] = 162'b111111111111111101000000000000001101111111111111111110000000000000000100000000000000000010000000000000000111000000000000001101000000000000000000000000000000010001;
    mem[148] = 162'b111111111111111110000000000000001100000000000000000100111111111111110110111111111111110011000000000000010011000000000000001010111111111111111011000000000000000001;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100111111111111111010111111111111111100;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule