`include "num_data.v"

module w_rom_25 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000011010000000000000001000010000000001000000001111111111101101011000000000011010101000000000100000010111111111100111010000000000000001101111111111111100101;
    mem[1] = 162'b000000000000011100111111111111101110000000001001011110000000000010100111000000000010100010000000000100101110111111111000100100000000000100101011000000001110001111;
    mem[2] = 162'b111111111110101011111111111110010100111111111101010111000000000000101101111111111111100000111111111101101001000000000000000000000000000000011000111111111011001101;
    mem[3] = 162'b000000001000110101000000011110100111111111111010111001111111100101001011000000010010001100111111101001011000111111110110111100111111110101001100000000000111101101;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111000001101111111111100000111111111111101100101000000000111100011111111111010111111111111111110010010111111111111100001111111111010111000111111111100001011;
    mem[33] = 162'b000000000100011101111111111100010111111111111111111010111111111101010000000000000000101110111111111110011100111111111011110110111111111100100101111111111111111100;
    mem[34] = 162'b000000000100100101000000000001111000111111111000101111000000000100000111111111111111001011000000000001100111000000000011011001111111111110110000000000001011010000;
    mem[35] = 162'b000000000010001110111111111010110111111111111110101011111111111011010111000000000010011101000000000100100000000000001100011000111111111011011110000000000101001011;
    mem[36] = 162'b000000000011100101000000000110100100111111111111110111111111110110101101000000000111010010000000000100001010111111111111001000000000000000010010000000001000110001;
    mem[37] = 162'b000000000010001111111111111100100000000000000110110111111111111000001111000000000000011100000000000111011111000000000100111001111111111101011011111111111101100100;
    mem[38] = 162'b111111111110010101000000000011100101000000000011111101000000000100000010000000001001010111000000000001101001000000000001100000000000000100100000000000000001110000;
    mem[39] = 162'b111111110111111001111111111110000101111111111011100001000000001001001011111111111101111100111111111100001010111111111110011010111111111100000111111111111101101100;
    mem[40] = 162'b000000000100011011000000000000101111000000000001010101111111111010011110000000000001000111000000000100101001000000000011110111000000000011100111111111111110111101;
    mem[41] = 162'b111111110001101011000000001001110001000000000000000000111111111011001100000000000101000000000000000101001010000000000010111100000000000110100010111111111101000001;
    mem[42] = 162'b000000000010011111111111111111110101111111111101100011111111110011101101000000000010011010000000001000110000111111110110011110000000000010011100000000000000010110;
    mem[43] = 162'b111111111100101011000000000011011011000000001000010101111111111000110001000000001010011101000000000101100011111111111111111100000000001010000001000000000110011110;
    mem[44] = 162'b000000000100010110000000000010110001111111111111111011000000000100111110111111111011110111111111111100101001111111111011100010111111111000001001000000000011101111;
    mem[45] = 162'b111111111010011011111111111111001100000000001001001110000000000100101110111111111110110111000000000000011111000000000000110111111111110110110111000000001001001000;
    mem[46] = 162'b111111111011001110000000000101011010111111111111011010111111111110000011000000000001000100000000000000000100111111111000100000000000000101110100111111111001100110;
    mem[47] = 162'b000000000011110101000000000101001001111111111010011100000000000011111100111111111010100110000000000000110011111111111001000111000000000110110110000000000000111110;
    mem[48] = 162'b111111111011101011111111111101000001000000000000001010111111111111001101111111111111101100111111111101010100000000000000100101000000000100011111111111111110010100;
    mem[49] = 162'b111111111010010011111111111001010001000000000010110111000000000000100100111111111100111001000000000011100101111111111100100001111111111101100001111111111100010011;
    mem[50] = 162'b000000000000011001000000000010111101111111111001100010000000000100111001111111111110001011000000001000000001000000000011000011000000000110111000111111111011011001;
    mem[51] = 162'b000000000010000000000000000011011000000000000001001011000000000100001010000000000011111101000000000001011001000000000011001000000000000011101001111111111100011110;
    mem[52] = 162'b000000001000000010000000000110110110000000000100100101000000000011101001111111111111010101000000000111010100000000000001011110000000000011011011000000000000111101;
    mem[53] = 162'b111111111110000111000000000010010100111111110101110001000000001000111010000000000100011000000000000001011101111111110110110011111111111011011101000000001001001100;
    mem[54] = 162'b111111111011001111111111111111101100111111111010001100000000000101000010111111111100001101000000000100100000000000000001111001111111111011001100111111111111001101;
    mem[55] = 162'b111111111110011001111111111011110100000000000011101101000000000110011100111111111111110010000000000110000011000000000100011111000000000110000111111111110110001001;
    mem[56] = 162'b111111111101001111111111111111010101111111111110001000111111111111000101111111111101110011000000000010101010000000000011101000111111111111010001111111111011001000;
    mem[57] = 162'b000000000000000001111111111100010111000000000011010011000000000001000101111111110111101001111111111111111100111111111011001100111111111110000010111111111011001100;
    mem[58] = 162'b111111111100101101000000000011000010111111111110000001000000001001001111111111111111001110000000000100100000000000000000000010111111111101001001000000000011000110;
    mem[59] = 162'b000000000010011110111111111101110000000000000011111111000000000010100101111111111100011011111111111111010110000000001101101011111111110010000001111111110001011011;
    mem[60] = 162'b000000000010101111000000000001111000111111111101111011000000000010101101111111111111101010111111111111000100000000000001111101111111110110010001000000000100110000;
    mem[61] = 162'b111111111010111111000000000010100110111111111110110011000000000111111011000000001000100011111111111111010110111111111001111111000000000111100101111111111100010001;
    mem[62] = 162'b111111111110100111000000000111000000111111111111110110111111111111100100111111111111100011111111110111000011000000000101100110000000000000111011000000000010010110;
    mem[63] = 162'b000000000001011110111111111101111111000000000011101111000000000110010010000000000010111101111111111101110110111111111111011000000000000011110110111111111111001001;
    mem[64] = 162'b000000000100000100000000000010101011000000000001110011000000000001110011111111111011110101000000000100100111000000000010000111000000000011111010000000000001011000;
    mem[65] = 162'b000000000011110010000000000111111100000000001001100010000000000011110000000000000000110010111111111111000100000000000010011011000000000010000000000000000000000110;
    mem[66] = 162'b000000000100100111000000000010110000000000000110001110000000000011100100111111111011011100111111111101010111000000000101001011111111111000001001111111111011101001;
    mem[67] = 162'b000000000110101010000000000100010011000000000011111011000000000101110100000000000001100000111111111110001011000000000100000001111111111101011010111111111101010001;
    mem[68] = 162'b000000000000010110000000000101010000000000000010111010000000000000111010111111111100011010111111111110100001000000000101001100000000000000111001000000000011011011;
    mem[69] = 162'b000000000101000101000000001000110110000000000110010011000000000011001111111111111110110010111111111110000110111111111111111101111111111100111101000000000000010100;
    mem[70] = 162'b000000000110010001000000000100001011000000001001110001000000000010111000111111111100101010111111111110011001000000000101101110111111111110011011000000000001101001;
    mem[71] = 162'b000000001001110110000000000110101110000000000000100111000000000100011110111111111101110100000000000011110011000000001000001111111111111111011011000000000000011000;
    mem[72] = 162'b000000000010101110000000000100000110000000000011000100000000000011101001000000000010110100111111111000111110000000000010101110111111111011000111111111111100101101;
    mem[73] = 162'b000000000000100111111111110111100000111111111010110001111111111010111100111111111010100110111111111010101111000000000011111110000000000011011111111111111100100100;
    mem[74] = 162'b000000000011100000000000000001110010000000000101001110000000000010101101111111111110100100111111111011110011000000000100011111111111111011101101111111111100110001;
    mem[75] = 162'b000000001100110010000000001101111100000000010010100011000000000110000001000000000011000001000000000101111100000000000101001100000000000011001011000000000101010000;
    mem[76] = 162'b000000000111010000000000010001001000000000010001110110000000001000001101000000000111101011000000000100100101000000001010100000000000000011100001000000001001111100;
    mem[77] = 162'b000000001011111001000000001101111011000000001100111001000000000111101010000000000010110111111111111111100010000000000110001111111111111111001111111111111111110101;
    mem[78] = 162'b000000010000000100000000010001011001000000010011001110000000001011101110000000001001011000000000000111111010000000001011000110000000000001111011000000000101010010;
    mem[79] = 162'b000000001001100101000000001000011111000000001010111000000000000011110111000000000000100101000000000000100100000000000011010001111111111100010110000000000010111010;
    mem[80] = 162'b000000000110110010000000000001101000000000000111010000000000000101000001000000000100101010111111111111010111000000000010110011111111111101110000000000000000001110;
    mem[81] = 162'b000000000101010101000000000010101000000000000010111010000000000010100110111111111101010010000000000011000001000000000010111111111111111110011010111111111111111101;
    mem[82] = 162'b000000001001111010000000001010010000000000001010001100000000000111011101000000000100101101000000000010100101000000000011010000000000000001001010000000000001001011;
    mem[83] = 162'b000000001011011011000000010001100101000000010001011000000000000111001110000000000000011101000000000010111111000000000110000001000000000000000101000000000010000111;
    mem[84] = 162'b000000000011000011000000000110111100000000000011101001111111111011011101111111111011000000000000000110001100000000000000000000111111111110100100000000000011000100;
    mem[85] = 162'b000000000110001110000000000110101110000000001100101111000000000111010100000000000011000000000000000100001011000000000101101111000000000000101100000000000101111110;
    mem[86] = 162'b000000001110000000000000010000001011000000010000111110000000001100010010000000000110100111000000000100100111000000001100011001000000000101110100000000001110011011;
    mem[87] = 162'b000000000110111001000000000011010111000000000101101100000000000101001000000000000100101110111111111100010110000000000100110010000000000011110000000000000001101011;
    mem[88] = 162'b000000000011100010000000000111001010000000000100011001000000000001100010111111111110110100111111111111101100000000000010110111000000000000001001111111111011000101;
    mem[89] = 162'b000000000100010101000000001010110010000000001011101010111111111110011100111111111111111111000000000010011001000000000010100000111111111110001110000000000011111110;
    mem[90] = 162'b000000000110001101000000001110000001000000001001011110000000000101111110000000000000111100000000000000111010000000000111100100000000000100001001000000000010111011;
    mem[91] = 162'b000000000011101011000000000011111110000000001000111100000000000011011100000000000011010111000000000000110011000000000100101011000000000000101110000000000100111110;
    mem[92] = 162'b000000000001010000000000001000010000000000000111111100000000000110011111000000000000100110000000000010110101000000000011101000000000000001001111111111111101011011;
    mem[93] = 162'b111111111100111000000000000010001101000000000011001100000000000000000101111111111010000100000000000000100010000000000001000100111111111100110101000000000000110010;
    mem[94] = 162'b000000000001000000000000000011110000000000000010100110111111111100100100111111111010100111111111111100100100000000000010110011111111111111011110111111111010000010;
    mem[95] = 162'b000000000011100111000000000111111010000000001010101100000000000100011011111111111101010001000000000011110100000000000010000010000000000000001101000000001000001010;
    mem[96] = 162'b111111111000111011111111111011110111000000000000010101000000000000001011000000000000001001111111111110111101111111111111100101000000000000001000111111111110110110;
    mem[97] = 162'b000000000000010011000000000000000010000000000010010011111111111111001110000000000000010010111111111111001000000000000000001101111111111111010110111111111111100010;
    mem[98] = 162'b111111111101010100000000000000111101000000000010101110000000000000010011000000000000001111111111111111110000000000000000001100111111111110111101000000000000111101;
    mem[99] = 162'b111111111111110010111111111000010000000000000010010001000000000001000101111111111111101111111111111111101000111111111010010111111111111111100001000000000000010001;
    mem[100] = 162'b000000000000011010000000000111100101000000001101100000111111111010011110111111111101101100000000000011101001000000000000100100111111111111000001111111111111101111;
    mem[101] = 162'b000000000000100110000000000001111110000000000011001111000000000000101010111111111111110011111111111111011011111111111110001000111111111111011101000000000000000101;
    mem[102] = 162'b111111111000111110111111111101110111000000000011000010111111111110100101111111111111010010000000000000110100000000000001111000111111111011111011000000000000110001;
    mem[103] = 162'b111111111111110010000000000000000101000000000001010010000000000000001100111111111111000010111111111101101110000000000010000010000000000001111011111111111011110100;
    mem[104] = 162'b111111111010000101111111111110000010000000000001011100111111111111001001111111111111111011000000000000000111111111111111110110111111111111100101111111111110001000;
    mem[105] = 162'b000000000000100001000000000000000000000000000010010110000000000001000011000000000000001101111111111110100101000000000010010001111111111001101010111111111100101111;
    mem[106] = 162'b000000000000001111000000000000001111111111111111110011111111111111011001000000000000111100111111111110001000111111111001001110111111111101110110111111111111110100;
    mem[107] = 162'b111111111101110010111111110111010110111111111010111010111111111010000101111111101101010000111111110001101101111111111110111110000000000000111011111111111111011101;
    mem[108] = 162'b000000000000000001000000000000111101000000000110011101111111111111100101000000000000001010111111111111011110000000000001001100111111111111000101111111111110110110;
    mem[109] = 162'b111111111111111010111111111101011111000000000101001111111111111101111111111111111110101011000000000001110010000000000010101110111111111011101001111111111011110110;
    mem[110] = 162'b111111111011010000111111111111111101000000000100001101111111111111111001000000000000011110111111111100100101111111111101011111000000000000010001111111111110100000;
    mem[111] = 162'b111111111001110100111111111111110001000000000101000111000000000000000100111111111111101110111111111111111000000000000001011111000000000000001000111111111110000100;
    mem[112] = 162'b000000001100110010000000001001111001000000011011101010000000000011101110000000000010010000000000000100110011000000000101001111000000000101000110000000000001101000;
    mem[113] = 162'b111111111111101100111111111110110100000000000110100100111111111110111001111111111111100010111111111111011001000000000000110011000000000001011010111111111110110101;
    mem[114] = 162'b000000000000011010000000000000111100000000001011110011111111111101010100111111111111101100000000000000001101111111111110001110111111111010110000111111111011001110;
    mem[115] = 162'b111111111110011001111111111111001101000000000110000101000000000000110110111111111001001110111111111110110100000000000010001101111111111110100011111111111111111111;
    mem[116] = 162'b111111111111100010000000000001100011000000000000000111111111111111110100111111111111010010000000000001000001111111111111100100111111111111111101111111111110011101;
    mem[117] = 162'b111111111110100111111111111110100011000000000011011000111111111100010010111111111110011111111111111011110011000000000000100101000000000000000100111111111110101010;
    mem[118] = 162'b111111111101111100111111111101010010000000000010100010111111111111100000000000000000011111111111111110101101111111111111110100111111111100110101000000000001011001;
    mem[119] = 162'b111111111110100111000000000000010001000000000001100011111111111101110100000000000000100101111111111111100101111111111111000100111111110111110111111111111010100101;
    mem[120] = 162'b111111111101111010111111111111111110000000000001011110000000000000100110111111111110110101000000000000101101000000000001011110111111111111111010111111111111000111;
    mem[121] = 162'b000000001001111001000000001000000000000000010110010101000000000001110110000000000000100001000000000011111111000000000011011110000000000110100111000000001000010111;
    mem[122] = 162'b000000000000011011111111111100011010111111111111011110000000000000011000111111111111111110111111111110110010000000000000100011111111111111110011111111111110111001;
    mem[123] = 162'b111111111111000110000000000000001001000000000000011110000000000000011001111111111111111010000000000000001001000000000000001001111111111111110001111111111011101010;
    mem[124] = 162'b111111111110110010111111111110011110000000000010101000111111111111010010000000000000001011111111111110111111111111111110001101111111111101100111111111110100001010;
    mem[125] = 162'b111111111101011011111111111100010010111111111100110110111111110010010001000000000000001111000000000000000011000000000000110001111111111110111111000000000000000000;
    mem[126] = 162'b111111111111110100000000000000001100000000000001010000111111111110101010000000000000110011111111111111001010000000000000010001000000000000010000111111111101110111;
    mem[127] = 162'b000000000000100001000000000000011100000000000000011001000000000000001110111111111110100000000000000000010100111111111111110111000000000000100011000000000000100100;
    mem[128] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[129] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[130] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[131] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[132] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[133] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[134] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[135] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[136] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[137] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[138] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[139] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[140] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[141] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[142] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[143] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[144] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[145] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[146] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[147] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[148] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule