`include "num_data.v"

module w_rom_15 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000110111110111111110110110000111111111101110111000000000011011010111111110111011011111111111110000011111111111111001010111111111011110100000000000001111110;
    mem[1] = 162'b000000000000101110111111111010010111111111110110000110000000000001101110111111110111111101000000000000001011000000000010001111111111111100010001111111111111100111;
    mem[2] = 162'b111111111101010010000000000001010110000000000001101001111111111111001101000000000101011100111111111111001100111111111011001011000000000001010000000000000011000101;
    mem[3] = 162'b000000010100000110111111110001000100111111101101010101000000000101010101111111110111011100111111110100101101000000000001000111000000001011010110111111110001100100;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b000000001000000110111111111101101100111111111101110001000000000010010001111111111010000001111111111110010011000000000111100101111111111001101000000000000000100110;
    mem[33] = 162'b111111111011110111000000000011011110111111111011001011000000000100101001111111110010111010111111111111101111111111111101110110000000000101100101111111111110011010;
    mem[34] = 162'b111111111111100111000000000101100101111111110111000101111111111011000001000000000000000010111111111001100010000000001010001010111111111000010111111111111011000000;
    mem[35] = 162'b111111111100101001000000000100101001111111111100111011000000000001011010111111111100001011000000000000000010111111111101100011000000000101100010111111111011010000;
    mem[36] = 162'b000000001000010010111111111010001000000000000010000010000000000000100001000000000010010100000000000101000010000000000000110101111111111011011011000000000011111111;
    mem[37] = 162'b111111111111001110111111111110010001000000000000000110111111111101110001111111111000100001111111111111111101111111111011101011000000000100010100111111111111100001;
    mem[38] = 162'b000000000010101010000000000011100011111111111111111110000000000110010011000000000010101100000000001001001010000000000101000101000000000100101101000000000100011011;
    mem[39] = 162'b000000000001010000111111111100011001000000000001101101111111111100101000000000000000010110000000000010000011000000000011001101111111111110100010000000000011111001;
    mem[40] = 162'b000000000001111100000000000101101101000000001001101100111111111110000100000000000010010010111111111110110100000000000100011001000000000111001001000000000001010111;
    mem[41] = 162'b111111111101010111000000000000100111111111111101100111111111111010100000111111111011110100111111111011000111000000000011001000111111111001010111000000001001001011;
    mem[42] = 162'b000000000010001000111111111101000111000000000011000101111111111100011011000000001000101101111111111000110011111111111101010010000000000100001101000000000010000110;
    mem[43] = 162'b000000000000110100111111110111000001000000000001000011111111111000110111111111111011110101111111111001111110111111111011001000000000000001111010111111111100000001;
    mem[44] = 162'b000000000100110111000000000001110010111111110111001110000000000011101010111111111101010101111111111000111001111111111100010101000000000000100101111111111110000111;
    mem[45] = 162'b000000000001011010000000000011100011000000000111101010111111111101010101111111111101110100000000000100101001111111110111000110000000000010000001000000000100110001;
    mem[46] = 162'b111111111111111100111111111100010101000000000100111101111111111101001101000000000010100001000000000010010101111111111001001110111111111001010000000000000101000001;
    mem[47] = 162'b111111111000111100000000000001000101000000000001011010111111111011000010000000000011011111111111111010111001111111111101101111111111111010111111111111111001100101;
    mem[48] = 162'b111111111100010111000000000011111000000000000001111111000000000010111111000000000111101110000000000001110101000000000100111001111111111010000011000000000100010111;
    mem[49] = 162'b000000000110111000111111110101111100111111111100000010000000000111001010000000000010000111111111111010100110111111110101010110111111111101111011111111111010001010;
    mem[50] = 162'b111111111101001100000000000010101111111111111001111100111111111111101010111111111110100001000000000011111000000000000010111000000000000101001101111111110111101111;
    mem[51] = 162'b000000000110011101000000000101010001000000001010001010000000000110011111000000001001101111000000001001011011000000000010111011000000000110111100000000000100110101;
    mem[52] = 162'b000000000000000000000000000000111001000000000011011000000000000111111011000000000011111100000000001000111000000000001011100110000000000001001101000000000010010000;
    mem[53] = 162'b111111111001110000000000000110000001111111111100000001111111111110010101111111111111110001111111111011001110000000000001111110000000000011111100000000000100100011;
    mem[54] = 162'b111111111111110011111111111011101101111111111110010011111111111111011010000000000110111011000000000000100101000000000010111110000000000100010110000000000000001000;
    mem[55] = 162'b000000000001111111111111111011110010111111111001101101111111111101000101111111111011000110111111111101001100111111111110010001111111111011010100111111111001011011;
    mem[56] = 162'b000000000001110011111111110101011100000000000100011011111111111101010001111111111111001111000000000111110011111111110111110010111111111111001011000000000101111000;
    mem[57] = 162'b000000000100010011000000000000110001111111111011111000000000000111011101111111111011111111111111111111111011111111110100111000000000000000010001111111111011111111;
    mem[58] = 162'b000000000001111001111111111111001100111111111111111100000000000010110010111111111011010011000000000101101001111111111111000111000000000001100010000000000010100001;
    mem[59] = 162'b000000000001110000000000000101011011111111110110000100000000000000111110000000000010110101000000000010111101111111110100111110111111111010011011000000000100011100;
    mem[60] = 162'b000000000000001011000000000110000110111111111100100011000000000010111110111111111101111110111111111000101010000000000011000110111111111111100001111111111110000111;
    mem[61] = 162'b111111111101001111111111111100000110000000000001010110000000000001110100000000000101111111111111111101001101000000000101101111111111111000110101111111111101011000;
    mem[62] = 162'b000000000010111000000000000101111000111111111111111000111111111110001100000000000100110100111111110101111110000000000100110011111111111100110010111111111011100010;
    mem[63] = 162'b111111111110011011000000000000101001000000000100010101000000000000111010111111111110000010000000000001010011000000000010110100111111111101001001000000000001000100;
    mem[64] = 162'b111111110110101001000000000000010100000000000001111100000000000011110101111111111101010000000000000011100000111111111110100100000000000010100011000000000001101100;
    mem[65] = 162'b000000000001000110111111111111010001111111111011100001000000000000001000111111111110011010000000000011001011111111111111010100000000000001001010111111111110100101;
    mem[66] = 162'b111111111110101111111111111010001001111111111001111000000000000000101101000000000100110001111111111000010010000000000011100110111111111100111111111111111001011000;
    mem[67] = 162'b111111111101011011111111111110000010111111111011101001000000000001110111111111111100111010000000000000010000111111111010100001000000000100011011111111111101001101;
    mem[68] = 162'b000000000000001000111111111111010011111111111100010110111111110111111110000000000001100101111111111101001100000000000000101101111111111011011111000000000101100011;
    mem[69] = 162'b111111111100101000000000000010101010000000000100110111111111111110011100000000000001010010111111111101110111000000000001111111111111111111100100000000000000010010;
    mem[70] = 162'b000000000011011110111111111111011001111111111100010001111111111000111000000000000001111111111111111110011110000000000000011110000000000100111001000000000100011010;
    mem[71] = 162'b111111111110001100111111111111110001111111111111000101000000000001001110000000000010011011111111111110110110000000000100001110111111111111011001000000000000100010;
    mem[72] = 162'b111111111100001110111111111101101000111111111101010001000000000001111111111111111101000000111111111011110100111111111011110000111111111101011110111111111110111001;
    mem[73] = 162'b111111111101001010111111111011100101111111111100000000000000000011101011000000000000011111000000000100110001000000000001111010111111111010011111000000000000010000;
    mem[74] = 162'b111111110111010010000000000100111110111111111100101110111111111101110001111111111101000001000000000000011000000000000010011110111111111010111110000000000001010001;
    mem[75] = 162'b000000000001011001000000000010100100000000000010010111111111111111001001111111111110011011111111111100110100111111111111110000111111111110100001111111111101101101;
    mem[76] = 162'b000000000111010110000000000001111011000000000100001000000000001000111100000000000101110011000000000001111010000000001000100100000000000010110001000000000100000000;
    mem[77] = 162'b111111111011111111000000000101011010111111111101001100000000000000100001111111111100010000111111111101101011111111111110011100111111111101011010111111111100001100;
    mem[78] = 162'b000000000000110110000000000101000100000000000010101010000000001100000101000000000001110100000000000010000111000000001010010000000000000010000000000000000010010011;
    mem[79] = 162'b000000000001001101111111111110110111000000000001101110000000000100001001000000000000010001111111111111110000111111111101111010000000000110000110111111111011111111;
    mem[80] = 162'b111111111100110101111111111101011101111111111010011100000000000010010011000000000011110001111111111101001000111111111101011011111111111111100010111111111110001001;
    mem[81] = 162'b000000000010001100111111111001000001111111111011001001000000000000010100111111111111110010000000000010111011111111111111101111111111110110000000000000000001010110;
    mem[82] = 162'b000000000001111000000000000000011100111111111100110110000000000010101011111111111001000111111111111111000111111111111011010100000000000010000001111111111100111111;
    mem[83] = 162'b000000000001010010000000000011100001000000000001111110000000000100010001000000000000110111111111111111100011000000000000100101000000000011001000000000000111011111;
    mem[84] = 162'b000000000010010101000000000010001000111111111100101111111111111111011111111111111111011101000000000001001111111111111010000111111111111100011110000000000001010111;
    mem[85] = 162'b000000000001110000000000000001001000111111111111100101000000000111010111111111111100010001000000000011000100000000000000010110000000000001011100111111111100101000;
    mem[86] = 162'b111111111100000111111111111110111100000000000010111111000000000111010110000000000100101110000000000011101000000000001000001100000000001000010111000000000011101011;
    mem[87] = 162'b111111111100111100111111111111110100000000000001011001111111111100011100111111111100110101111111111111010010000000000011000001111111111111110001000000000000100111;
    mem[88] = 162'b000000000010111010000000000000110110000000000000000100000000000010111010111111111001011100111111111100111010111111111101001100111111111111101100000000000011101010;
    mem[89] = 162'b111111111100001111111111111101110110111111111101100101111111111010010111000000000010001101000000000101010101111111111110001111000000000000101001111111111011111010;
    mem[90] = 162'b111111111100001101000000000010000101000000000110001011111111111111100001111111111111000110000000000010000100111111111010111011111111111110110001000000000010111011;
    mem[91] = 162'b111111111011110010000000000010101001111111111110010100000000000010011001000000000010001101111111111101100010111111111101010100000000000001111001000000000000000001;
    mem[92] = 162'b111111111010010001000000000000010011111111111111111011000000000001111100111111111110000101111111111011111010000000000000100111111111111010100110111111111100100001;
    mem[93] = 162'b111111111101111100111111111101101111111111111001111101111111111101001010000000000100011011111111111110011100000000000001101110111111111101001001000000000000111100;
    mem[94] = 162'b000000000010100110111111111110110001000000000011000011111111111010001101000000000010111000000000000001110010111111111100110010111111111100111111111111110111000010;
    mem[95] = 162'b000000000000110001111111111101000000111111111000110001111111111111110000111111111111011010000000000000101110000000000101101110111111111011101001000000000011000110;
    mem[96] = 162'b111111111111111111111111111111111001000000000000001011000000000000010000000000000000001101000000000000011100111111111111110011111111111111101101111111111111111100;
    mem[97] = 162'b000000000000000111000000000000001010000000000000000000000000000000011011000000000000000001111111111111111001000000000000000000111111111111110000000000000000010011;
    mem[98] = 162'b111111111111101101000000000000001110111111111111101101000000000000011100000000000000010000111111111111111110000000000000001110000000000000010010111111111111110000;
    mem[99] = 162'b000000000000011000000000000000011010000000000000000101000000000000000000000000000000001110000000000000001010111111111111101000111111111111111001111111111111101110;
    mem[100] = 162'b000000000000011000000000000000001001111111111111111101000000000000001101000000000000000111000000000000000110000000000000001011000000000000011100000000000000001100;
    mem[101] = 162'b000000000000000011000000000000010001000000000000011001000000000000001110111111111111111100111111111111110110111111111111100111000000000000001000000000000000010001;
    mem[102] = 162'b000000000000001110111111111111111001111111111111111010111111111111110101000000000000000010111111111111111011000000000000000110000000000000000000000000000000011001;
    mem[103] = 162'b000000000000001101000000000000011110000000000000000001000000000000001110000000000000010011000000000000000000000000000000001100111111111111111100111111111111101001;
    mem[104] = 162'b111111111111111000000000000000010110000000000000011000000000000000010101000000000000001001000000000000011100000000000000010011000000000000001111000000000000001011;
    mem[105] = 162'b000000000000001110111111111111111010000000000000001001000000000000010010111111111111110111111111111111110110000000000000000010111111111111101011111111111111100001;
    mem[106] = 162'b000000000000001111000000000000001110111111111111111011000000000000000101111111111111111111000000000000000110000000000000000101111111111111110101000000000000010010;
    mem[107] = 162'b111111111111110000111111111111110100111111111111111100111111111111110011111111111111111010111111111111111011000000000000010101000000000000100100000000000000010010;
    mem[108] = 162'b000000000000100000000000000000011010000000000000011010000000000000000000000000000000010101000000000000001101000000000000010100111111111111111100000000000000000110;
    mem[109] = 162'b000000000000001110000000000000010100000000000000000000000000000000010010000000000000000011111111111111111100111111111111111101000000000000000100111111111111111100;
    mem[110] = 162'b000000000000000110000000000000000100000000000000001101111111111111110101111111111111111111111111111111111010000000000000011100111111111111101110000000000000010100;
    mem[111] = 162'b000000000000000010000000000000000001000000000000010101111111111111111000000000000000001110000000000000000110000000000000000011000000000000000101000000000000011110;
    mem[112] = 162'b000000000000110001000000000000011111000000000000111010000000000000001110000000000000001011000000000000011111000000000010001010000000000000010010000000000000011001;
    mem[113] = 162'b000000000000000001111111111111110101000000000000011101000000000000000100000000000000001000000000000000000101111111111111110011111111111111111111000000000000011010;
    mem[114] = 162'b111111111111111110000000000000010101000000000000001111000000000000000010000000000000000011000000000000010001000000000000010000111111111111111101111111111111111110;
    mem[115] = 162'b111111111111111110111111111111110110111111111111111001000000000000010011000000000000010000000000000000001011000000000000010000000000000000001001000000000000010001;
    mem[116] = 162'b111111111111101010111111111111111011111111111111111000111111111111111001111111111111110111111111111111111010111111111111100110111111111111111101000000000000010100;
    mem[117] = 162'b000000000000001000111111111111111011111111111111111111000000000000010100111111111111111111000000000000000001000000000000001110111111111111111011000000000000000010;
    mem[118] = 162'b000000000000101000000000000000000001111111111111110110000000000000001110000000000000000010111111111111111110000000000000011011000000000000010000000000000000100000;
    mem[119] = 162'b000000000000010010000000000000010011000000000000000011000000000000001101000000000000001000000000000000001011000000000000001000000000000000001101000000000000011111;
    mem[120] = 162'b000000000000001000000000000000000000000000000000001100000000000000000011000000000000010001000000000000010111000000000000011000000000000000010011111111111111111110;
    mem[121] = 162'b000000000000100000000000000000010101000000000000100010000000000000011100000000000000001110000000000000101111111111111111000111000000000000100010000000000000110101;
    mem[122] = 162'b000000000000001100000000000000011011111111111111111000111111111111111011111111111111111000111111111111111101000000000000001000000000000000010001000000000000001001;
    mem[123] = 162'b000000000000001001000000000000011001000000000000010011111111111111110100000000000000000010111111111111111100000000000000000111111111111111111001111111111111110110;
    mem[124] = 162'b000000000000001110000000000000010001000000000000010010000000000000000010111111111111111001000000000000001001111111111111110110111111111111111111111111111111111000;
    mem[125] = 162'b111111111111101010111111111111101111111111111111101111111111111111111110111111111111110100111111111111111110000000000000010011000000000000000001000000000000001011;
    mem[126] = 162'b000000000000000010000000000000010100111111111111101011111111111111101110000000000000000011000000000000010101111111111111111001000000000000000010000000000000001110;
    mem[127] = 162'b111111111111101010111111111111111100000000000000011011111111111111110000111111111111101110111111111111100111111111111111111001111111111111110001111111111111111100;
    mem[128] = 162'b111111111111111110000000000100000101000000000110111000000000000011111100111111111100000001111111111111110011000000000000100110111111111111101110000000000001101111;
    mem[129] = 162'b111111111111111100111111111111111001000000000000000000000000000000000000111111111111111110111111111111111111111111111111101000000000000000000001111111111110101011;
    mem[130] = 162'b000000000000000010000000000000000000000000000000000011111111111111111011000000000000000001111111111111111100000000000000000011111111111111110100111111111111111011;
    mem[131] = 162'b000000000000000101000000000000000001111111111111110111111111111111111000000000000000000000111111111111110100111111111111111100111111111111110111111111111111111010;
    mem[132] = 162'b111111111110101011000000000000010000000000000000001001111111111111100010111111111111111110111111111111001001000000000000010000000000000000010101000000000000101101;
    mem[133] = 162'b111111111111110011111111111111111010111111111111111001111111111111111111000000000000001000111111111111111101000000000000110101111111111111111110000000000010011011;
    mem[134] = 162'b000000000011001101000000000101001000000000000101001001111111111111111100000000000000000111111111111111111010111111111111111101111111111111111111111111111111110101;
    mem[135] = 162'b000000000000010000111111111111111001111111111110010010111111111111111101111111111110010101000000000011011111000000000000000101111111111111010011000000000101001101;
    mem[136] = 162'b000000000000000111111111111111111011111111111111110001111111111111111010111111111111111100111111111111111000111111111111111100000000000000001000000000000000000000;
    mem[137] = 162'b111111111111110101111111111111110111111111111111110000000000000000001011000000000000000001111111111111111101111111111111111100000000000000000000000000000000001010;
    mem[138] = 162'b000000000000000011000000000000000000000000000000000011111111111111111010000000000000000001111111111111110100111111111111110110000000000000001110000000000000001000;
    mem[139] = 162'b111111111111111011111111111111111101000000000000000001111111111111111110111111111111111111111111111111111001000000000000000011000000000000000100111111111111111101;
    mem[140] = 162'b000000000010100101000000000011010101000000000101101100000000000010010010111111111111101110000000000000101111111111111111010011000000000000011001111111111100111111;
    mem[141] = 162'b111111111111110101111111111111111111111111111111111010000000000000000111000000000000000001111111111111111111000000000011011110000000000011000000000000000001011010;
    mem[142] = 162'b000000000101100111000000000101000110000000000011110100111111111111110000111111111111110111111111111111110101111111111111110100000000000000000000111111111111111111;
    mem[143] = 162'b000000000011011111111111111110111111111111111111100101000000000000101000000000000000111110000000000000110010111111111111110000111111111111101001000000000100000101;
    mem[144] = 162'b111111111111111110000000000000000010000000000000000011111111111111111110111111111111111111111111111111111111000000000000000101000000000000000010000000000000000010;
    mem[145] = 162'b111111111111111111000000000000000011111111111111110111000000000000000111000000000000000010000000000000000011000000000000000000111111111111111110000000000000000001;
    mem[146] = 162'b000000000000000111000000000000000010000000000000000001000000000000000100000000000000000011000000000000001011000000000000001110000000000000001000000000000000000010;
    mem[147] = 162'b111111111111111010000000000000001000000000000000000101000000000000000000000000000000001110111111111111111110111111111111111010111111111111111000000000000000000010;
    mem[148] = 162'b111111111111110101111111111111111111111111111111101100111111111111110010111111111111101011111111111111111110000000000000001011000000000000000011000000000000000000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110111111111111111110111111111111111001;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule