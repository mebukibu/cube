`include "num_data.v"

module w_rom_3 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000001101111000000000001110000111111110100010011000000000001000100000000000101000011000000000110001011111111111110001000111111111111100010111111111100111001;
    mem[1] = 162'b111111111100111110000000001100101000000000001001101011000000001001111011111111111110011100000000001101010100111111111101111000000000000100100001000000001001100001;
    mem[2] = 162'b111111111110001011000000000000010011111111111100111011111111111011101000000000000010111110111111110001100110111111111110111101111111111111111110000000000100110111;
    mem[3] = 162'b111111110100110010111111101010011100000000011000000011111111110111010001000000000011111000000000001101111110111111111011111001111111110111010010000000001011001001;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b000000000000001100000000000000110111000000000100011001000000000110010110000000000011101010111111111110011100000000000101100000111111111010001010111111111101111011;
    mem[33] = 162'b000000000001010011111111111111101111111111111000101010111111111000011001000000000000000011000000000110011110000000000101011111000000000001101110111111111101101100;
    mem[34] = 162'b000000000110000001111111111111100100111111111111100100000000000000110001000000000000010100111111111101000111000000000111010111000000001100101111111111111101011101;
    mem[35] = 162'b000000001001010110000000000000001010111111110100010010000000001000011101111111111111111000111111111101101001000000000101100010000000000000000010111111111111000011;
    mem[36] = 162'b111111111110010010000000000011111111000000001001100011000000000001000001000000000000010100000000000001100000000000000111001101000000000000110111000000001101100011;
    mem[37] = 162'b111111111011010011000000000001001011000000000100001101111111111101110111000000000100100110000000000011110000000000000100100101111111111110000010000000000000010100;
    mem[38] = 162'b000000000011110010000000000011010010000000000000011001000000000000000000000000000011101111000000001001001101000000000100111100111111111011111010000000001010000100;
    mem[39] = 162'b111111111100010110000000000111001100111111111010000011111111111101110110111111111111010000111111111001010010111111111011111001000000000000110101000000000001011111;
    mem[40] = 162'b000000000001101000000000000001100010000000000010101011111111111110100000000000000011010011111111111110010011111111111001000101000000000000101100000000000101100010;
    mem[41] = 162'b111111110101111001111111111110111010000000000000111001000000000101100001000000000001101101111111111111101000000000001000010001111111111100101110111111111110111000;
    mem[42] = 162'b000000000111101000000000000100010110111111111101011111111111110111101010000000000100111111000000000100101101111111111101100011000000000010110110000000000100101000;
    mem[43] = 162'b000000000001010101111111110101110110000000000101001101000000000010000101000000000110100000000000000011100110111111111111101100000000000100100100000000000101110110;
    mem[44] = 162'b000000000000010101111111111111110101111111111010001010000000001010110111000000000010000100111111111010101011111111111010010010000000001000011001111111111101111000;
    mem[45] = 162'b000000000010110001111111111010010010000000000000000111111111111011111000111111111011100001000000000000111110000000000010111011111111110100111111000000000100000100;
    mem[46] = 162'b000000000011000100111111111001001001111111111100101111111111111110000111111111111111110011111111111100010111000000000001000111111111111111011111111111111100001100;
    mem[47] = 162'b000000000100110100111111111001101011111111111111010100000000000001011000000000000110111001111111111011110100111111111101101011000000000010010110111111111011000001;
    mem[48] = 162'b111111111100101110000000000001111010000000000110110101111111111100011000000000000000110001111111110001110111000000001000101011111111111011010001111111111110111010;
    mem[49] = 162'b111111111111101011000000000010000010000000000000100110000000000001101011111111111100111000111111111010001110111111111100011101111111111110001000111111111110110110;
    mem[50] = 162'b000000000101111011000000000110100001111111111101101001111111111001110111111111111101110001111111110101110011000000000110001100000000000100100011000000000011100111;
    mem[51] = 162'b000000001000010001000000000100110001000000000100101001000000000100001010000000000011000010000000001001010000000000000110110100000000000010110001000000001011010111;
    mem[52] = 162'b000000000101110111000000000000001100000000000010110101000000000010011101000000000001111001000000001001000110000000000011000111000000000101000000111111111100110111;
    mem[53] = 162'b111111111110010101111111111100100111111111111100011010111111111100101100111111111011100000111111111111011111000000000001101010000000001000100110000000000000001001;
    mem[54] = 162'b111111111111000001000000000100110100000000000101111110111111111001100110000000000111011011111111111111100010000000000010011100111111110111111110111111111101001000;
    mem[55] = 162'b000000000101111001000000001001010100111111111000010110111111111110011000000000000010110101111111111000101100111111111111100000111111111111100111000000000011110101;
    mem[56] = 162'b111111111011001000111111111111010000000000000001110011000000000000101000111111111100010101111111111100100001000000000000001000111111111010010100000000001001101111;
    mem[57] = 162'b111111111100101100000000000100011111000000000011010101000000000100000101111111110111011001111111111111010111111111111010111100000000000100111001000000000010010001;
    mem[58] = 162'b000000000001010011000000000110111001111111111110011100111111111000011100000000000010001110000000001000101010111111111111001110111111111000011010000000000010110101;
    mem[59] = 162'b111111111001111001111111111100110100000000000100111110000000000101101011111111110111111111000000000101110001000000000010101101000000000001001100111111110100100110;
    mem[60] = 162'b111111111111110100000000000110010010111111110111000101000000000010110100111111111101100110000000000011111010111111110110101001000000000111110000111111111100100101;
    mem[61] = 162'b111111111101011110111111111101101110111111111101010000111111111101000010111111111101010010000000000010001010000000000010001000000000000100011011111111110110100101;
    mem[62] = 162'b000000000110011110111111111111011111111111111111001001000000001010001110111111111110000101000000000010001100111111111110100100000000000111100000000000000000001001;
    mem[63] = 162'b000000000100100000000000000000110100000000000010011001111111111101000101000000000110001010000000000000100101111111111101000001000000000110101100111111111010100011;
    mem[64] = 162'b111111111011100101111111111101001010111111110101001110111111111110000001111111111011111001000000000000110001000000000000011100111111111111011000111111111011111101;
    mem[65] = 162'b111111111111011110111111111011100011000000000100001101000000000000011101000000000100101100111111111100111101000000000010000110000000000011111010000000000000001110;
    mem[66] = 162'b000000000100000000000000000010000100000000000000011001111111111110001100111111111100001111111111111100111101111111111111110100000000000001111100111111111100011000;
    mem[67] = 162'b111111111101001001111111111001110101111111111110110010111111111110101101111111111010011000111111111111001101000000000101100010111111111110001110000000000001001010;
    mem[68] = 162'b111111111101101011111111111011100100111111111001010000000000000000101000000000000001101110000000000000101100111111111100001001111111111110101101111111111110100011;
    mem[69] = 162'b000000000001110111000000000011110010111111111111011100111111110101011110111111111101001100111111111110110010000000000001101011000000000100001001000000000000111010;
    mem[70] = 162'b000000000001111111000000000010000100111111111101111110111111111011011011000000001001011110111111111111010100111111111001110110000000000100010011000000000100010010;
    mem[71] = 162'b000000000101010000000000000010110000111111111101101000000000000000100011111111111110001111111111110100101101111111111110001001000000000000101101111111111100001100;
    mem[72] = 162'b111111111011001101000000000000010011111111111111111101111111111111111101111111111110101101000000000000111001111111111111010111000000000110110001111111111100000100;
    mem[73] = 162'b111111110110110111111111111111010011111111111111010010111111111010001111000000000010111101000000000001101001000000001001010101000000000101000101111111111001111100;
    mem[74] = 162'b111111110101101100111111111111111100000000000010100000000000000001000110000000000101111111000000000000110000111111111111000010111111111100000101111111111101010110;
    mem[75] = 162'b000000001001001100000000001011110001000000000101100011000000000001010011000000000000110001111111111011010011111111111111000100111111111011111001111111111100111101;
    mem[76] = 162'b000000000100110100000000000100010000000000000111001100000000000100111111000000000000010010000000000000110011000000001011000100000000001010101111000000001001111000;
    mem[77] = 162'b000000000000100001111111110110101110000000000000101110000000000000100110000000000001000110000000000000100011000000000001111011111111110111001101000000000000010100;
    mem[78] = 162'b000000001000101011000000001001110011000000000100011101000000000101100001000000000110110111000000000000100100000000000001100100000000000010000100000000001010001101;
    mem[79] = 162'b000000000001101100000000000001101000000000001010111010000000000010000011000000000001000010111111111011010011111111111111001000000000000000111101111111111101000101;
    mem[80] = 162'b111111111111010010000000000000001000111111111010010111000000000011100011111111111010100011111111111101010101111111111100000010111111111011100111000000000010010111;
    mem[81] = 162'b111111111100110111111111111101011101111111110110000000111111111110110110000000000010010100000000000000100010111111111001000110000000000001011101111111111101111111;
    mem[82] = 162'b000000000000100110000000000001001100000000000000000001000000000101010111000000000000111010000000000110101111111111111011011110111111111100100110000000000010101110;
    mem[83] = 162'b000000001000100001111111111111101111000000000000001011000000000000010100000000000011100000000000000001101100000000000000110110000000000000101111000000000011110011;
    mem[84] = 162'b111111111101101000111111111111111101111111111111111111111111110010011111111111111110000010111111111111111011111111111100101000000000000010101111111111111111101001;
    mem[85] = 162'b000000000011110111000000000010001001000000000011100000000000000011011011111111111111111001000000000010111001111111111101110000000000000011100010000000000101110110;
    mem[86] = 162'b000000000010110111000000000011111100000000000011111001000000000010101101000000000110101000111111111011111001000000001001010001000000001010101110000000001001001110;
    mem[87] = 162'b111111111100111011111111111010110110111111111111000101111111111110010101111111110111110011111111110100000001111111111110010100000000000000011001111111111111001111;
    mem[88] = 162'b000000000001100101000000000001011100111111111011100011111111111100100101111111111111000101111111111101000001111111111101010110000000000000111111000000000101101110;
    mem[89] = 162'b111111111100101010111111111101011100000000000100010011111111111010010110111111111111011101111111110101111000111111111101101010111111111011011000000000000011111110;
    mem[90] = 162'b111111111111001000000000000010100011111111111110101011111111111101001111000000000101010101111111111100110010111111111011010101000000000000000111111111111101000111;
    mem[91] = 162'b111111111111101001111111110110100010111111111000010011000000000001100000000000000011101100111111111100001101000000000110000001000000001010010000000000000010000100;
    mem[92] = 162'b000000000001010011111111111011010000111111111011100001000000000001111011111111111111001011000000000100000100111111111000000111111111111101000111000000000000101010;
    mem[93] = 162'b111111111111011101111111111110000001000000000001101101111111111011111111111111111111100111111111111011101100111111111100111010111111111101101101000000000001110110;
    mem[94] = 162'b000000000010100011111111111110000001000000000000100000000000000011100100000000000000011001111111111110100011000000000010101001111111111100101010111111111101010101;
    mem[95] = 162'b000000000001111001000000000000110000000000000010111000000000000011001011111111111100011000000000000011101100111111111110110110000000000011101011000000000010100110;
    mem[96] = 162'b111111111111111000000000000010101110111111111100001000111111111110001011111111111110110111000000000010011111000000000001110101111111111111101110111111111100011000;
    mem[97] = 162'b111111111110111010000000000001011001111111111100111011000000000010100010111111111100111101111111111011111100000000000101000111000000000100110011111111111101111001;
    mem[98] = 162'b000000000011101000000000000000010011111111111101101001111111111110000111000000000010111100111111111101101001000000000100101010111111111111001010111111111101100010;
    mem[99] = 162'b111111111101001000000000000010101001000000000001011001111111111111101001111111111110100110111111111001000000000000000010101111000000000001111000000000000001100000;
    mem[100] = 162'b000000000011110001000000000001101000000000000011010011000000000010111001000000000001001110000000000001111011000000000010111111000000000100111111000000000000001011;
    mem[101] = 162'b111111111111000110111111111110101001111111111111111001111111111101001001111111111101101001000000000001010011000000000001011001000000000010100011111111111110001011;
    mem[102] = 162'b111111111110000101111111111111011101111111111110001000111111111110100011111111111101001010000000000010001001000000000101110110000000000011011000111111111111111001;
    mem[103] = 162'b000000000000101101111111111101001101111111111111111101000000000000101110111111111000110110000000000001010001000000000011110111000000000000010000111111111111111000;
    mem[104] = 162'b111111111111110111111111111111110000111111111101010011111111111110111000111111111100000101111111111110000110000000000011001101000000000111101110000000000010000011;
    mem[105] = 162'b000000000010001100111111111111110110000000000010110000111111111010001110111111111111001000111111111111111110000000000000110010111111111100001100111111111010010101;
    mem[106] = 162'b111111111110100110111111111110100001111111111110001000111111111111110111111111111101001010111111111101001101000000000100101001000000000001001001111111111011101100;
    mem[107] = 162'b111111111011010001111111111111111001000000000010010010111111110111101110111111111111111000111111111001011001000000000011100010111111111110110111111111111111011111;
    mem[108] = 162'b111111111101000100111111111110010000000000000000010111111111111110001110111111111111100101000000000100101011000000000101110001111111111001011010111111111110011011;
    mem[109] = 162'b111111111011100111111111111110100110000000000001110010111111111010010010111111111010011100111111111100101100111111111111111000111111111011011000111111111100110001;
    mem[110] = 162'b111111111101111001000000000001011101111111111111101111111111111101101010111111111110111111000000000000100011000000000011001000000000000001000100111111111110101100;
    mem[111] = 162'b000000000000110111111111111100100101111111111111110111000000000010011100111111111111000001000000000010001001111111111111001100000000000011010101000000000010000011;
    mem[112] = 162'b000000001000101001000000000111000110000000000111000000000000010000001110000000001000011101000000000011101011000000011111100011000000001101101001000000000111100101;
    mem[113] = 162'b000000000011000100111111111101011011000000000000001110000000000000001010000000000000111010000000000000101001000000000011110101000000000001001000000000000001001110;
    mem[114] = 162'b000000000000000000000000000001100101111111111110000110000000000000110001111111111101001101000000000000100000111111111110100111111111111101110110111111111101111010;
    mem[115] = 162'b000000000000011101111111111111110111000000000001001010111111111101010100111111111111100100000000000010000101000000000101001101111111111101001101111111111111100010;
    mem[116] = 162'b000000000010010100111111111011100011111111111110100011111111111100000100111111111111101110000000000001011011000000000011011011000000000001101001000000000010100011;
    mem[117] = 162'b111111111111110110000000000001010001111111111110111101111111111101010101111111111111110000111111111100010010000000000011110001000000000001111101111111111110000010;
    mem[118] = 162'b000000000001101000000000000001111010000000000000000011000000000000111011000000000000101011111111111111111100000000000001100000111111111110001101000000000000101100;
    mem[119] = 162'b111111111101011010111111111110010010111111111101011100111111111110101100111111111110000111000000000000100000000000000001000001111111111110111101111111111101010100;
    mem[120] = 162'b111111111111010000000000000001010100000000000000100011000000000000101100000000000001010110111111111100100100000000000011101001000000000010101111111111111100111100;
    mem[121] = 162'b000000000111001110000000000100001010000000000100011010000000001101010011000000001010001000000000000110101100000000101000010101000000010100110010000000001100010100;
    mem[122] = 162'b111111111111100100111111111100010100000000000100010001000000000010100010111111111011010000111111111100110100000000000110100100111111111110110011111111111111111101;
    mem[123] = 162'b000000000100010110111111111111100011111111111111001010111111111101100100000000000000010110111111111110000101000000000000100000000000000001101011000000000001010011;
    mem[124] = 162'b111111111001100000111111111110101000111111111101010001000000000000011111111111111110000110000000000000010101000000000001100111000000000001001110000000000100101011;
    mem[125] = 162'b111111111011001111111111111001110110111111110101111101111111111110101111000000000000000000111111111111101101000000000010101010000000000001100100000000000000100101;
    mem[126] = 162'b111111111110100011111111111110010110000000000000110100000000000000111111111111111111011011000000000010011110000000000101011101000000000001010001000000000000000101;
    mem[127] = 162'b000000000001011010111111111111011001000000000000011001000000000000000010000000000000111101000000000000010111000000000100011111111111111111010110000000000010000011;
    mem[128] = 162'b111111111111000111111111111111111110111111111110010101111111111111001110111111111110100111111111111111011101000000000010011100000000000001110111111111111110110110;
    mem[129] = 162'b000000000000000011111111111111111110000000000000000011111111111111111110111111111111111100000000000000000110000000000010000100111111111110111110111111111110111111;
    mem[130] = 162'b111111111111111110111111111111110101111111111111111111000000000000001000000000000000001110000000000000010001000000000000010000000000000000000001000000000000000010;
    mem[131] = 162'b000000000000000011000000000000001000000000000000010001000000000000001011111111111111111100000000000000000101000000000000001100000000000000000010000000000000000000;
    mem[132] = 162'b000000000100110111000000000010100110000000000000000011000000000101101011000000000101001101000000000000000100000000000000001001111111111111101110111111111111100111;
    mem[133] = 162'b111111111111111101111111111111110111000000000000000010000000000000000100111111111111111100000000000000000001000000000000010001000000000011101010000000000011010110;
    mem[134] = 162'b111111111111111010000000000000000001000000000000001101111111111111111001000000000000001001000000000000000010111111111111111101111111111111111110111111111111111000;
    mem[135] = 162'b111111111110111011111111111111100101111111111111110000111111111111011101000000000010010000000000000011100010111111111111010001000000000000000101000000000000111000;
    mem[136] = 162'b111111111111011000111111111111101001000000000001000100111111111111110001000000000001010110111111111111111111000000000001100010000000000000001011000000000001011011;
    mem[137] = 162'b000000000000000000000000000000000000000000000000000001000000000000000110111111111111111101000000000000000111000000000010110000000000000101001110000000000011001010;
    mem[138] = 162'b111111111111101001000000000000111000111111111111100000000000000000001100000000000000000110000000000000000111000000000000000110000000000000000000000000000000001011;
    mem[139] = 162'b000000000000100000000000000000011100111111111110111011111111111111111001000000000000000001111111111111110101000000000000100111111111111111101100000000000001010101;
    mem[140] = 162'b000000000000001000000000000000010100000000000000000111000000000000001100000000000000010110000000000000000001000000000000000100111111111111111011111111111111111100;
    mem[141] = 162'b111111111111111110000000000000000011111111111111110101111111111111111111111111111111111010111111111111111110111111111111111110111111111111111111000000000000000111;
    mem[142] = 162'b000000000000001000111111111111111110111111111111111100111111111111111101111111111111110111000000000000000111000000000000000101111111111111111101111111111111111011;
    mem[143] = 162'b000000000000001010000000000000000011000000000000000100000000000000000010000000000000000010000000000000000011000000000000000000111111111111111100111111111111111110;
    mem[144] = 162'b000000000000000001111111111111111110000000000000000110000000000000000000000000000000000100111111111111111101111111111111111110111111111111111100111111111111111010;
    mem[145] = 162'b111111111111111000111111111111110110000000000000000010000000000000000000111111111111111101000000000000000111111111111111111110000000000000001001000000000000000110;
    mem[146] = 162'b000000000000001011111111111111111110000000000000000000111111111111111101111111111111110110111111111111111011000000000000000101111111111111110111111111111111110010;
    mem[147] = 162'b111111111111111010111111111111111101111111111111110011111111111111110110111111111111111110111111111111111010111111111111111001000000000000000010000000000000000111;
    mem[148] = 162'b111111111111111100000000000000000010111111111111110111111111111111110011111111111111110010000000000000001000000000000000000100000000000000001001111111111111111001;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000111111111111111010000000000000000010;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule