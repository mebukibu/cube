`include "num_data.v"

module w_rom_30 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b111111111110011001000000000111010010000000000010101100000000001000001011000000000101001001000000000100011110111111111000101100111111111111100100111111111110101111;
    mem[1] = 162'b000000001011110110111111111011101101111111110101000010111111111100000011111111101110110001111111110000101011000000000100010000000000001011000110111111101110010001;
    mem[2] = 162'b111111111111101010000000000011000111111111111101011011111111111010101001111111111110010001111111111111111100111111111011001010000000000101010010111111110110111110;
    mem[3] = 162'b000000001101100001000000001000100001111111101111100001000000001110001111111111111111111010111111111001010010000000000100010001111111111111001100111111101101011001;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111100101010111111111111110010111111111111011100000000000010010101111111111001111000000000000101001110111111110110000011111111110110001001111111111110111101;
    mem[33] = 162'b111111111101111011000000000000010001000000000100010101000000000010110011111111111110001100111111110101101101000000000101101011000000000110000111111111111101001100;
    mem[34] = 162'b000000000000101100111111111010010001000000000001101011000000001010010101000000000000100001000000000001100111000000000010100010111111111110100101000000000000001010;
    mem[35] = 162'b000000000111000010111111111001001111000000000101100100111111111110101001111111111101100101000000000111111111000000000111011000111111111110100010111111111100011010;
    mem[36] = 162'b111111111110011010000000000101001011000000000001010101111111111010110101000000000010111001111111111101111000111111111000101100000000000011010101000000000001011001;
    mem[37] = 162'b000000000000010010000000000010001111111111111110011100111111111100100101000000000001001011111111111101001100000000001000010100111111111010011000111111111110110010;
    mem[38] = 162'b000000000010001111000000000110101000111111111100100010000000000100000101000000001000110101000000000110010001000000000011101101000000000011111001111111111011101010;
    mem[39] = 162'b000000000101101100000000000000000101111111111110100101000000001001001011000000000101101010000000000101110011111111110110110011000000000000001101111111111011001011;
    mem[40] = 162'b111111111110111110000000000111111001000000000100110001111111111111110010111111111110000111111111111011000110000000000000000011000000000111010001000000000010000111;
    mem[41] = 162'b111111111101011010111111111110011010111111111101100110111111111101001010111111111100100100111111111010100001000000000010101111000000000110010101000000000110011110;
    mem[42] = 162'b111111110111111101111111111001100000111111111111111000000000000011010111000000000011010101000000000110100101111111111010011000000000001000111101000000000100011111;
    mem[43] = 162'b000000000001000110000000000111110000000000000111000100111111111000011110000000000110010100111111111101101000111111111000010010000000000101000011111111111011111001;
    mem[44] = 162'b000000000001110100000000000001100100111111111010101101000000001001111111111111111101100111111111111001001000000000000011001000111111111111011100111111110011110100;
    mem[45] = 162'b111111111111010100111111111101001001111111111011100000111111111111010100000000000011000111111111111101110010000000000011110011111111111111101110000000000000001100;
    mem[46] = 162'b111111111110001000000000001000100100111111111101011100111111111101001010000000000100000101111111111000101000111111111101001110000000000101011100111111111000100101;
    mem[47] = 162'b000000001001011010111111111010000001111111111110101101111111111110000001111111111001010100000000000001000010111111110111110101000000000011011011000000000001011101;
    mem[48] = 162'b000000000001100110111111111101000110111111110110101100111111111101001011000000000000100001000000001010100011000000000100101101111111111110010011111111111110000011;
    mem[49] = 162'b111111111101001011000000000010001100000000000000000110111111110111101000000000000000111101111111111000100111000000000111000100000000000001000111111111111101100110;
    mem[50] = 162'b111111111101000001111111111110011101111111111001000100111111111111011011000000000101000111111111110111111110111111111100000100000000000010101010000000000001011000;
    mem[51] = 162'b000000000001000111000000000010000101000000000110011010000000000010110011000000000111110110000000000001011101000000001000000111000000000011101101111111111100010101;
    mem[52] = 162'b111111111110001111000000000100000100111111111111110000000000000001000111000000000011100100111111111101111101000000000001010100000000000101100101111111111111100001;
    mem[53] = 162'b000000000000100101000000000101001011111111111110010111000000000000110110000000000010000010000000000001101010000000000001100110000000000011000001000000001001100100;
    mem[54] = 162'b000000000101010100111111111110101101111111110111010010000000000010010001111111111011101110000000000001111111000000000110100010000000000000010000000000000001110100;
    mem[55] = 162'b000000000011101001111111111010101010000000000100111001111111110110100000111111111101110111111111111110011100111111111110001110111111111001101001111111111110001000;
    mem[56] = 162'b000000000000010011000000000010100000111111111101010000111111111011101111000000000001001111000000000011111000111111111111001100000000000000010101000000001001011110;
    mem[57] = 162'b111111111101000001111111111110100001111111111011010011000000000101110100111111111100001110000000000100011010111111111111001010000000001000010010111111111100101011;
    mem[58] = 162'b000000000111001000000000000000011001000000000001011111000000000000101001000000000110101010000000000011010010000000000001000000000000000010011111000000000000011011;
    mem[59] = 162'b111111111011100101000000001000000101000000000001010011111111111011110111000000000010001011000000000110011101111111111111011100111111111111111100000000000000100110;
    mem[60] = 162'b111111111011100000111111111100010110000000000110001110111111111010110100000000000111110101111111111010000010111111111101110011000000000011110101111111111010011000;
    mem[61] = 162'b111111111100000000000000000110011100111111111101011010111111111010100100111111111111011000000000000111110011111111111110011101000000000011011110111111111111110111;
    mem[62] = 162'b000000000110000110000000000000111101111111111011110111111111111111000011111111111111011000000000000101101010111111110110110100111111111011101101111111110111010100;
    mem[63] = 162'b000000000110010100000000000010110101111111111010011010111111111110010111000000000001101001000000000000000010000000000111000010000000000101000000111111111000010000;
    mem[64] = 162'b111111111011010110111111111100100111111111111010110110111111111110010010111111111101011001000000000101011101000000000000011111111111111101101100111111111101111011;
    mem[65] = 162'b111111111101110001111111111100111011000000000001000011111111111101100001111111111010000111000000000010110111000000000010001001000000000011010011000000000010001001;
    mem[66] = 162'b111111111010000000000000000000101110000000000100000110000000000001111110111111111100010000111111111001001110000000000000000011111111111110011111000000000010000110;
    mem[67] = 162'b111111111011100001000000000100001110000000000100101011111111111111110111111111111111111101000000000000111111111111111100111011111111111100011011111111111011100110;
    mem[68] = 162'b111111111101000110111111111111100101000000000001111101111111111001001111111111111111111001000000000000011110111111111111011101000000000001010010111111111000111011;
    mem[69] = 162'b000000000000100001000000000001110011111111111111001001111111111011111011111111111111010011000000000101100111111111111110011101111111111100101001000000000101101110;
    mem[70] = 162'b000000000110001000111111111010101110111111111110011100000000000000000111111111111101010110000000000010111010000000000001000001111111111001110100111111111111010010;
    mem[71] = 162'b000000000100001000111111111111000010111111111111001111111111111110010010111111111100010101111111111101011101111111111110101101000000000000011010000000000000011011;
    mem[72] = 162'b000000000110001100000000000010110111111111111111011010111111111111001100111111111010111000111111111001001011111111111111100110000000000000001000111111110111011110;
    mem[73] = 162'b000000000001011101000000000001011011000000000011010010111111111111100111000000000000011100111111111110111001000000000110001110000000000010010111000000000001010111;
    mem[74] = 162'b111111111001111001111111111100001100000000000011010111111111111100001100111111111000001101111111111011101101111111111111111110000000000000011000111111111010100000;
    mem[75] = 162'b000000000000101011111111111111101100000000000111110000111111111110010010000000000000001110000000000100000000000000000010110011111111110110001111111111111001100001;
    mem[76] = 162'b000000000011101000111111111111001010000000000110111000000000000111111000000000000010000111000000000110010000000000000111100101000000000001110001000000001001001011;
    mem[77] = 162'b111111111111111101000000000001011011000000000011111100000000000110001100000000000000110100111111111111101001000000000000111100111111111000101110000000000111011100;
    mem[78] = 162'b000000001000101011000000000101000010000000000100000000000000000100101010000000000100010010000000000101010011000000000111111110000000000101010010000000000101101100;
    mem[79] = 162'b000000000010110001111111111101110101111111111110101000000000000000110010000000000010111100111111111101111110111111111111100000000000000000101001111111111110001111;
    mem[80] = 162'b000000000010011010111111111111101001111111111011010000111111111000011011111111111111101010111111111011000110111111111111001010111111111001111011000000000101110111;
    mem[81] = 162'b111111111110100100111111111111111010111111111100101101111111111101100101111111111101100110111111111100110011000000000011001101000000000000011110000000000100001100;
    mem[82] = 162'b000000000001011010000000000011101111000000000000100110111111111110101010111111111100010011111111111110100110000000000011100001111111111001011100111111111110100110;
    mem[83] = 162'b000000000101001000111111111010011101000000000111100111000000000011001111000000000101000011000000000110001010111111111101010110111111111111011100000000000001101011;
    mem[84] = 162'b000000000011100000111111111100001101111111111001010101000000000100001111111111111100111101000000000010110001111111111010111101000000000010010110000000000001101000;
    mem[85] = 162'b000000000110010011000000000000101000111111111111000011000000000011011000000000000010100010000000000011011010000000000011001001111111111011100011000000000011011010;
    mem[86] = 162'b111111111111111000000000000010011000000000000011100111000000000110001001000000000000111010000000001001010011000000000110011100000000000010000100000000000110110101;
    mem[87] = 162'b000000000100010011111111111110101100111111111101101011111111111110101100000000000010010000111111111110110111000000000001100110000000000010011011111111111100001110;
    mem[88] = 162'b111111111110000000000000000000101001111111111110100111111111111111111001000000000010111110111111111110111001000000000010000000000000000001001010111111111111001101;
    mem[89] = 162'b111111111100110101111111111111010001000000000011000011111111111101110111111111111101110101111111111011010110000000000000111010111111111101100100111111111011010000;
    mem[90] = 162'b000000000001110001000000000010101101000000000010010011000000000100001010000000000100110101000000000001111101111111111101010001111111111111100111000000000011011011;
    mem[91] = 162'b000000000000000110000000000001000010000000000010001001000000000011010101000000000000010010000000000010010001000000000011110100000000000100001100000000000011010100;
    mem[92] = 162'b111111111110101101111111111111101001000000000100111000111111111101111101111111111010011100000000000010001011111111111010100110111111111101111011111111111101111111;
    mem[93] = 162'b000000000000101110000000000010010110000000000100000101000000000001011000000000000001111000111111111100110100000000000000001101111111111011011100000000000011011010;
    mem[94] = 162'b111111111010010010111111110111100100111111111111100001111111111111100010000000000001011101111111111100000100111111111011111110000000000000101100111111111111010101;
    mem[95] = 162'b000000000101000110000000000001011101000000000100111111111111111101010010111111111101111100000000000000011000000000000011101110000000000101011011111111111011111001;
    mem[96] = 162'b111111111111110100000000000000000011000000000000001001111111111111111110000000000000000001000000000000011010000000000000010000000000000000010110000000000000000010;
    mem[97] = 162'b111111111111111010111111111111111011000000000000010001111111111111111111000000000000000011111111111111110001000000000000001000111111111111111011111111111111110100;
    mem[98] = 162'b111111111111111000111111111111111101111111111111101111111111111111110100000000000000000110111111111111110111111111111111110110000000000000000110000000000000001001;
    mem[99] = 162'b000000000000000011000000000000001001111111111111111111111111111111111111000000000000001001000000000000001001111111111111111011000000000000001001000000000000000101;
    mem[100] = 162'b000000000000000100000000000000000101000000000000001111000000000000000111000000000000001111000000000000001100000000000000000100000000000000001001111111111111110010;
    mem[101] = 162'b000000000000011001111111111111111010111111111111111110000000000000000010000000000000000110111111111111111010111111111111110101111111111111111000111111111111111101;
    mem[102] = 162'b000000000000000100000000000000000011111111111111111010000000000000000111000000000000000111000000000000010000111111111111111010000000000000000001111111111111111101;
    mem[103] = 162'b111111111111111001000000000000001000000000000000001100111111111111111000000000000000000111000000000000000001111111111111111010000000000000001111111111111111111110;
    mem[104] = 162'b000000000000011010000000000000000111000000000000001101000000000000011011000000000000010010000000000000001111000000000000010001000000000000010000000000000000000011;
    mem[105] = 162'b111111111111110111000000000000000110000000000000001110000000000000000010000000000000000111000000000000000000000000000000010000000000000000001111111111111111110010;
    mem[106] = 162'b111111111111111111000000000000000110000000000000000001111111111111111100000000000000001010000000000000001111111111111111111001000000000000000001111111111111111001;
    mem[107] = 162'b111111111111110111000000000000000000111111111111111110111111111111111010000000000000000101111111111111110101111111111111111011000000000000000011000000000000000010;
    mem[108] = 162'b000000000000011011000000000000001110000000000000010000000000000000010100000000000000000010000000000000000110000000000000001100000000000000000100000000000000001100;
    mem[109] = 162'b000000000000001110000000000000000010000000000000000110000000000000011101000000000000000010111111111111101111000000000000010010000000000000000110000000000000000101;
    mem[110] = 162'b111111111111111110000000000000001111000000000000000101000000000000000111111111111111111001000000000000011000000000000000001100000000000000001100000000000000011111;
    mem[111] = 162'b111111111111110010111111111111101010111111111111111111111111111111110100000000000000010000000000000000000000000000000000000100000000000000001000000000000000010101;
    mem[112] = 162'b000000000000000110000000000000100010000000000000010110000000000000100111000000000000001000000000000000000010000000000001010000000000000000001110000000000000010010;
    mem[113] = 162'b000000000000010101000000000000001101000000000000001010111111111111110110000000000000000000000000000000010010111111111111111101111111111111111010000000000000001001;
    mem[114] = 162'b000000000000000011000000000000010011000000000000000010111111111111110111000000000000000010000000000000000111000000000000000001111111111111111110000000000000001000;
    mem[115] = 162'b111111111111111111111111111111110101000000000000001101000000000000001011000000000000001101000000000000000111000000000000110000111111111111111110111111111111110100;
    mem[116] = 162'b111111111111100110111111111111100111000000000000000001111111111111100110111111111111111001000000000000001111000000000000000000000000000000001100000000000000001011;
    mem[117] = 162'b111111111111111100111111111111111101000000000000000110000000000000000011111111111111110000111111111111111101000000000000011010000000000000010000111111111111111000;
    mem[118] = 162'b000000000000010101000000000000011101000000000000010100000000000000100101000000000000010000000000000000010011000000000000001000000000000000010111000000000000000110;
    mem[119] = 162'b111111111111110011111111111111111110000000000000011100000000000000000100000000000000000101111111111111111001000000000000000011000000000000010000111111111111111111;
    mem[120] = 162'b000000000000010110000000000000001101111111111111111010000000000000011110000000000000001010000000000000001110000000000000010010000000000000010001111111111111111100;
    mem[121] = 162'b000000000000000110000000000000001000000000000000010011000000000000000010000000000000001110000000000000001011111111111111100110000000000000010011000000000000100000;
    mem[122] = 162'b000000000000000111000000000000010000000000000000000011000000000000000101000000000000000111000000000000000011111111111111011101111111111111111101000000000000001001;
    mem[123] = 162'b000000000000010000000000000000001010111111111111110110000000000000001111000000000000001010111111111111110011000000000000000100111111111111111010111111111111101101;
    mem[124] = 162'b111111111111111010000000000000000110000000000000000000000000000000001100000000000000001011000000000000001100111111111111111110000000000000000010000000000000001100;
    mem[125] = 162'b111111111111111000000000000000000111111111111111110110000000000000000001000000000000001000000000000000000011111111111111101011111111111111101101111111111111110011;
    mem[126] = 162'b111111111111111110000000000000001111000000000000010111111111111111111100111111111111111111111111111111111111000000000000000000000000000000001001111111111111111111;
    mem[127] = 162'b111111111111111000000000000000000000000000000000001001111111111111100110111111111111110110000000000000001000111111111111111010000000000000000010000000000000000111;
    mem[128] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[129] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[130] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[131] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[132] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[133] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[134] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[135] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[136] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[137] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[138] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[139] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[140] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[141] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[142] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[143] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[144] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[145] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[146] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[147] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[148] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule