`include "num_data.v"

module w_rom_22 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000001100111000000000101111010000000000011111100000000000010101111111111111001100110111111111100101111111111111111010110111111111011101000111111111100100000;
    mem[1] = 162'b111111111001000101000000001110111001111111111010001111111111111011100001000000000100111000000000001111010010111111110010100000111111110110111111111111110110000101;
    mem[2] = 162'b000000000010001000111111111110001010111111111101000010111111111101101110111111111110010011111111111110100000000000000001011101000000000110000011000000000000101101;
    mem[3] = 162'b000000001111010011000000001010110101111111110101101101111111110011101111111111111101000111000000001111101111000000000111111101111111110001100011000000000010000001;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111111010011000000000000110100111111111000111011111111111101011011111111111011100101111111111000101110111111111110001110111111110101011101111111110001011110;
    mem[33] = 162'b111111111110110000000000000110010111111111111110000110000000000110010011111111111100000010000000000001111100111111110111001011000000000011110110111111111110011111;
    mem[34] = 162'b111111111010000110000000000001111110111111110111001010111111111100111000111111110111110010000000000000010001111111111110111111111111111010101011111111111010100000;
    mem[35] = 162'b000000000100101010111111111100101000111111111111010111111111111010011110111111110001110111000000000010111000111111110101111001000000000001110001000000000010000111;
    mem[36] = 162'b000000001011000001000000000011101010000000000010110001000000000011110001000000000100010110000000000110111010000000000000010010111111110111101010111111110010001111;
    mem[37] = 162'b111111111111000101111111111111111000000000001000000011000000000110000110111111110111111101000000000001010001111111111100000010111111111100100001000000001000101100;
    mem[38] = 162'b000000010110000010000000001000010001000000000100111011000000000011110010000000000101001101000000000111011011000000000110011000000000000001100010000000000010011011;
    mem[39] = 162'b000000000011111011000000000011111000111111111110000110111111110101101111111111111111101000000000000001110001000000000001000001000000000010111001111111111100111001;
    mem[40] = 162'b000000010110111100000000001010000011000000010000011010000000000011001101000000000000000101000000001000111111111111111111001111000000000101101101111111111110001101;
    mem[41] = 162'b000000001001111101111111111000010111000000001101011010111111110110100111111111111010111111000000000001100111111111111111111011111111111111100001111111111111001101;
    mem[42] = 162'b000000001001110101000000000110101111000000001000111110000000000010100101000000000100001001000000000000100111000000000010110010111111111100110001111111111101000011;
    mem[43] = 162'b000000000101001001000000000011100101000000000001110100000000000110101000000000000010000000000000000101000111111111111110110001111111110101101000000000000000101110;
    mem[44] = 162'b000000001010010010000000000100011110111111111101101010000000000001110011000000000101100001111111111010110100000000000011010010000000000111001000111111111001100010;
    mem[45] = 162'b000000001101110111000000000000100010000000000110010010111111111101000001111111111100111010000000001101101000111111111101011110000000000000010011111111111011100001;
    mem[46] = 162'b000000000100001100000000000010110011000000000001110011111111111100100111000000001001101001111111111111100010111111111111100001000000000010101100111111110110111101;
    mem[47] = 162'b000000000010100000111111111101010111111111111100100010111111111100111110000000000110110011111111111010011101111111111101010110000000000011001000111111110101011001;
    mem[48] = 162'b000000000001000110111111111100110011000000000000001100111111111111001000000000000010010101000000000000010011000000000001011101111111110110010001111111111000010100;
    mem[49] = 162'b111111111110100111111111111100100001000000000000110010111111111101110000111111111110001101000000000110011011000000000111001100000000000101001110000000001001010011;
    mem[50] = 162'b000000000100101011000000001000100000000000000100111100000000000101100011000000000100111010111111111111010110111111111101111001111111111110011000111111111111111000;
    mem[51] = 162'b000000100011100011000000001101011000000000001110101000000000001000011101000000001001101011000000001101001011000000000101010011000000000000000001000000001000111110;
    mem[52] = 162'b000000011000100001000000001110011000000000001000000010000000000100101100000000000101110101000000000101011011000000000011000100111111111110110000111111111100110111;
    mem[53] = 162'b000000000100010001111111111111110100000000000000000100000000001000101100111111111010010001111111111011011011111111110111100111111111111011010011000000000011000111;
    mem[54] = 162'b111111111101101110111111111011111000111111111100011111111111111000011011111111111110001101000000000001110100000000000100101000111111110011110111111111111100100111;
    mem[55] = 162'b000000000000100111000000000101100001000000000100001100000000000101101001111111111001101111111111111011000100111111111110111001000000000101101011000000000000101011;
    mem[56] = 162'b000000000011110011111111111010101101000000001000110111111111111011010011111111111001101010000000000000100001000000001001111101111111111001010100111111111101010010;
    mem[57] = 162'b000000000001011011000000000011010110111111110101101111000000001001000000111111111000100101111111111100110001000000000011111111111111111110111011000000000000010110;
    mem[58] = 162'b000000001011010011000000001000101000000000000100100101000000000000110110000000000001111101000000000011000000000000000100110110111111111000011011111111111011110111;
    mem[59] = 162'b000000001000000110111111111101000100111111111111101101000000000000101011111111111111101100111111110101111001000000000000000100000000000000111010000000000101001111;
    mem[60] = 162'b000000001011001110000000000010100100111111111011101111000000000000100001111111111001110110000000000000100000111111111100110100000000000000001110111111111110111110;
    mem[61] = 162'b000000000010110011000000000101101010111111111000010011111111111110010000000000000011010011000000000110011101111111111100001111000000000000101110000000000010010011;
    mem[62] = 162'b000000001110011100000000000011110001000000000001000100000000000010100110111111111010111101000000000100101101000000000100100000111111111110110110000000000011101000;
    mem[63] = 162'b000000001001111100000000001100000000000000000110000001000000000011001001000000000001110011111111111101100110000000000100100001111111111100010111000000000000110010;
    mem[64] = 162'b000000000000011101111111111110111101111111111010100001000000000011100011000000000001000110000000000000010100111111111111000001000000000011100000000000000000011011;
    mem[65] = 162'b111111111101000001111111111101000010000000000001010010111111111011110000000000000000111011111111111010011101000000000001100000000000000101010100111111111011000110;
    mem[66] = 162'b000000000001000110111111111110011010000000000011000011111111110110110110111111111010011110111111111111100100000000000110000101000000000000000011000000000001110001;
    mem[67] = 162'b111111111101101001111111111111111010000000000010001010000000000100110001111111111001001011000000000011101010111111110111110001111111111010110011111111111110000110;
    mem[68] = 162'b111111111100101000000000000010111111000000000101100110111111111100111111111111111001000100000000000011100100111111111101010111111111111011000011111111110011000011;
    mem[69] = 162'b111111111111111110000000000011010010000000000110011100111111111001110011111111111011011001000000000000111111000000000000110100111111111100101100000000001000110101;
    mem[70] = 162'b111111111111001110111111111100010011000000000110010011000000000101001110111111111111111110000000000100010100000000000010111110111111111001101101000000000101111110;
    mem[71] = 162'b000000000010011111111111111011000010000000000101000011000000000011010001111111111101110001111111111101101100111111111101010000111111111111010110000000000000010100;
    mem[72] = 162'b000000000001110101000000000011000100111111111011111011000000000101011110111111111100011101111111110101111101111111111101101001000000000011000010111111111100100100;
    mem[73] = 162'b111111111001100000111111111100010010000000000000010000111111111100110100111111111101101110111111111100001110111111111110111001000000000000101110111111111101110100;
    mem[74] = 162'b000000000101011001111111111010001100000000000110011010111111111011101010111111111010011110000000000001001101111111111000001000000000000011010000111111111100100101;
    mem[75] = 162'b000000000000011011000000000101111011000000000110110101000000000011011100111111111100001100111111111101010010111111111110011100111111111110010110111111111110001111;
    mem[76] = 162'b000000000001000110000000000110000011000000000100110111000000000001011010000000000001111100000000000001110100000000000011010101000000000101000010000000000100101001;
    mem[77] = 162'b000000000000010011000000000010010010000000000110101110000000000001101000000000000001110100000000000011110100111111111110110111111111111010111010111111111010010000;
    mem[78] = 162'b000000000100110110111111111111101111000000000101111000000000000100100100000000000101101101000000001000000110000000000001100111111111111111111011000000000010101111;
    mem[79] = 162'b000000000000001001000000000110001011111111111111111011000000000010001001000000000001000001000000000101011000000000000001011001000000000000000101111111111111111111;
    mem[80] = 162'b111111111000101010111111111110110101111111111111011011000000000000101110000000000110101111000000000010100011111111111001110111000000000000000110000000000111110100;
    mem[81] = 162'b000000000000011101000000000010010011000000000010001000111111111110100000000000000100100110111111111011110110111111111100010001000000000010010111111111111100101101;
    mem[82] = 162'b000000000001100111111111111100000000111111111110011010000000000110000001000000000101011010000000000011010110111111111010111000111111111101111000000000000010110111;
    mem[83] = 162'b000000000001101110111111111100110110000000001000011110000000001000000111000000000100100000000000000001110100111111111110011100111111111101111101000000000000100010;
    mem[84] = 162'b111111111100101011111111111110011110000000000001110010000000000000001111000000000010010110111111111110101001111111111110101101111111111011110100000000000011011100;
    mem[85] = 162'b000000000001100111000000000010110011111111111000011001000000000011001010111111111100111100000000000001000010000000000000100001000000001000000000000000000000011011;
    mem[86] = 162'b111111111100111010000000000001011111111111111011001101000000000001101011000000000001001001000000000101011111000000000101000100000000000100011011000000000110000111;
    mem[87] = 162'b000000000011101111111111111100101001000000000000110111111111111111001111000000000000100011111111111111110000111111111010000111000000000011000101111111111010101001;
    mem[88] = 162'b111111111110101000111111111111101011000000000010001011000000000100101111000000000011111000111111110110101000000000000101010011000000000010101011111111111110101111;
    mem[89] = 162'b000000000010100010111111111101111000111111111100101101000000000010001111111111111011010101000000000101000000111111111100000110111111111100110011000000000001011100;
    mem[90] = 162'b000000000001111000111111111111010100000000000111111011000000000010001100111111111111100000000000000110101101000000000101100100111111111101111010111111111101000110;
    mem[91] = 162'b000000000001000110000000000001010100000000000000100000111111111001110110111111111100001000111111111001101110000000000110000111000000000111101101000000000100010101;
    mem[92] = 162'b000000000011000011111111111110110101000000000100001111000000000001011011000000000000010101111111111101001011000000000001010101111111111001010110000000000111010011;
    mem[93] = 162'b000000000110111010000000000000010100000000000010101011111111111100100101000000000010110001000000000011000001111111111111001011000000000011000110000000000001100111;
    mem[94] = 162'b111111111010101011000000000011100001111111111111001010111111111110111101111111111011011010111111111100110100000000000000010000000000000101101001000000000111100101;
    mem[95] = 162'b000000000000101111111111111111110111111111111110011110000000000100010100000000000010100111000000000000110111111111111110011010111111111111000110000000000001100011;
    mem[96] = 162'b111111111111111010111111111111101001111111111111111010000000000000001000000000000000000001000000000000000100111111111111101011111111111111100101111111111111110011;
    mem[97] = 162'b000000000000000111111111111111110110000000000000000010000000000000001011000000000000000001111111111111111010000000000000000110111111111111110001111111111111111111;
    mem[98] = 162'b111111111111100101000000000000001101111111111111110111000000000000000111000000000000010000000000000000010001111111111111110100111111111111111110111111111111110001;
    mem[99] = 162'b000000000000011000000000000000010100000000000000011000000000000000000101000000000000001000000000000000000100111111111111111010000000000000000010000000000000000000;
    mem[100] = 162'b000000000000001111111111111111110011111111111111111001000000000000000010000000000000001010000000000000000000111111111111111010000000000000001111000000000000001000;
    mem[101] = 162'b000000000000001010000000000000011100000000000000100001000000000000000101111111111111111110111111111111110111111111111111100101111111111111111111000000000000010101;
    mem[102] = 162'b111111111111111001111111111111111010000000000000000010111111111111110100111111111111111111000000000000001111000000000000000101000000000000000101111111111111111100;
    mem[103] = 162'b111111111111111110000000000000010100000000000000000000111111111111111001000000000000001011000000000000000001000000000000000100000000000000000101111111111111110110;
    mem[104] = 162'b111111111111101110000000000000000010111111111111110101000000000000001001000000000000001011111111111111111111000000000000001010000000000000001010000000000000001111;
    mem[105] = 162'b111111111111110101111111111111110101111111111111101101000000000000001111000000000000000011111111111111111001111111111111111101111111111111110100111111111111111110;
    mem[106] = 162'b111111111111111101000000000000000000000000000000000111000000000000001000111111111111111111000000000000000110111111111111101110000000000000000100111111111111111000;
    mem[107] = 162'b111111111111111100111111111111111001000000000000000010000000000000000100000000000000000110000000000000000011000000000000000001000000000000001010000000000000000010;
    mem[108] = 162'b111111111111111010111111111111110101111111111111101100111111111111111100000000000000000101000000000000010011111111111111111110000000000000001000111111111111111101;
    mem[109] = 162'b000000000000010011000000000000000110000000000000001001111111111111111011000000000000000011000000000000001001000000000000010011111111111111111001111111111111111011;
    mem[110] = 162'b111111111111110110000000000000000111000000000000000101000000000000001000000000000000000100000000000000001001000000000000000111111111111111111011111111111111111001;
    mem[111] = 162'b000000000000010110000000000000000101000000000000001101000000000000001111000000000000001110000000000000001110111111111111110010111111111111111001000000000000001010;
    mem[112] = 162'b000000000000010110000000000000001101000000000000001001000000000000010000000000000000000100000000000000010001000000000000000001000000000000000000000000000000100000;
    mem[113] = 162'b000000000000001100111111111111110001000000000000000000000000000000001001111111111111111111000000000000000011000000000000001000000000000000001010000000000000000011;
    mem[114] = 162'b111111111111111110111111111111111000000000000000011110000000000000000000000000000000000001000000000000000111000000000000010010000000000000001111111111111111111100;
    mem[115] = 162'b111111111111111110000000000000001000111111111111110110111111111111110111111111111111111111111111111111110001000000000000001000000000000000000011111111111111111111;
    mem[116] = 162'b111111111111101110000000000000001000111111111111111100000000000000000100111111111111111110000000000000010111000000000000001000000000000000000100000000000000000111;
    mem[117] = 162'b000000000000000111111111111111111000111111111111000111000000000000010011111111111111110010000000000000000010000000000000010111000000000000000110111111111111111101;
    mem[118] = 162'b000000000000000111000000000000000011111111111111110011111111111111110010111111111111111000111111111111111011111111111111111010111111111111111100000000000000000101;
    mem[119] = 162'b000000000000001001000000000000011000000000000000011100000000000000000011000000000000001011111111111111110110000000000000000010000000000000001110000000000000000100;
    mem[120] = 162'b000000000000010000111111111111111111000000000000010011000000000000010110000000000000001111000000000000011010000000000000001001111111111111111010111111111111111110;
    mem[121] = 162'b000000000000000011000000000000001010000000000000001110000000000000001111111111111111111011111111111111111101000000000000110100000000000000001101000000000000100100;
    mem[122] = 162'b000000000000011101000000000000011000000000000000000100000000000000001011000000000000000000111111111111111100000000000000011011000000000000000110000000000000001111;
    mem[123] = 162'b111111111111110111111111111111101111000000000000010011111111111111111101111111111111110000111111111111110011000000000000001010000000000000000011000000000000000010;
    mem[124] = 162'b000000000000010001000000000000001000000000000000000011111111111111110111111111111111111100000000000000000001000000000000000110111111111111111010111111111111111001;
    mem[125] = 162'b111111111111111010111111111111110111111111111111100110000000000000000101000000000000001000111111111111111100111111111111110111111111111111111110111111111111110100;
    mem[126] = 162'b111111111111111110111111111111110011000000000000001100111111111111101110000000000000010110000000000000011010111111111111111000111111111111111001000000000000010111;
    mem[127] = 162'b111111111111110100111111111111111001111111111111101101000000000000000110111111111111101011111111111111100111111111111111111111000000000000000001111111111111111000;
    mem[128] = 162'b000000000000111010000000000100010001000000000100100101000000000101010100000000000001101000111111111111010111000000000010111101111111111111110101000000000000010111;
    mem[129] = 162'b111111111111111100111111111111111111111111111111111110000000000000000011111111111111111011111111111111110110000000000000100111111111111111011110000000000000000010;
    mem[130] = 162'b000000000000000010000000000000000000111111111111110011111111111111111110000000000000001000000000000000001011000000000000000111111111111111111101111111111111111100;
    mem[131] = 162'b000000000000001000000000000000000111000000000000000011000000000000000011111111111111111010111111111111110011111111111111111010111111111111110111000000000000001011;
    mem[132] = 162'b000000000001100001000000000001000111111111111110111001111111111111001111111111111111111000111111111111010100111111111111110010111111111111110010000000000000001010;
    mem[133] = 162'b111111111111111011111111111111111000000000000000000001000000000000000100111111111111110110000000000000000101000000000001100110111111111111111100111111111111101011;
    mem[134] = 162'b000000000110001111000000000011011000000000000101001000000000000000000111000000000000000111000000000000000100000000000000000000000000000000000000111111111111111100;
    mem[135] = 162'b111111111111111111000000000000101010000000000000000001111111111111110111000000000001100100000000000000111101000000000001000101000000000000011010000000000010111100;
    mem[136] = 162'b111111111111111110000000000000000100111111111111111111111111111111111111111111111111111110000000000000000101000000000000000100111111111111110111111111111111111110;
    mem[137] = 162'b000000000000000100111111111111111011000000000000000100111111111111111011111111111111111110000000000000001001000000000000000110000000000000001110000000000000000110;
    mem[138] = 162'b111111111111111000000000000000000010000000000000000011000000000000000101000000000000001111000000000000000000000000000000000000000000000000001010111111111111111110;
    mem[139] = 162'b000000000000010010000000000000001010000000000000001010000000000000000100000000000000001000000000000000000010111111111111111000000000000000000000000000000000000100;
    mem[140] = 162'b000000000100001100000000000000001000000000000010010100000000000001101100000000000001011101000000000000011110000000000001010001000000000001110001111111111100111010;
    mem[141] = 162'b111111111111110101111111111111111000000000000000000011000000000000000000111111111111110110000000000000000101000000000100010111000000000011011000111111111111100101;
    mem[142] = 162'b000000000100101010000000000010101011000000000010001111111111111111111010111111111111101101111111111111110001111111111111111000111111111111111000111111111111110101;
    mem[143] = 162'b111111111111101100000000000000001101000000000000001000111111111111111010000000000000000010000000000000101001000000000000000111111111111111101000000000000010010110;
    mem[144] = 162'b111111111111110100111111111111111000111111111111110100111111111111110011111111111111111100111111111111101101111111111111111001111111111111111101000000000000000001;
    mem[145] = 162'b000000000000000010111111111111111100111111111111111000000000000000000011111111111111101111111111111111110111111111111111110101111111111111100011111111111111101110;
    mem[146] = 162'b111111111111111101000000000000000011000000000000000011000000000000000000000000000000000011111111111111111101000000000000000011000000000000000011000000000000000101;
    mem[147] = 162'b000000000000001101000000000000000100111111111111111111111111111111111110000000000000000011111111111111111111111111111111111011111111111111111010000000000000000000;
    mem[148] = 162'b111111111111111110000000000000000101111111111111111011111111111111101111111111111111111001111111111111111000000000000000000010000000000000000001111111111111111110;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111101111111111111110101;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule