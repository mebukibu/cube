`include "../data/num_data.v"
`include "../data/state_layer_data.v"

module weight_store (
  input wire clk,
  input wire [2:0] cs,
  output reg valid,
  output reg [288*`data_len - 1:0] q
  );

  reg [10:0] addr;
  wire [`data_len - 1:0] ramout;

  reg init;
  reg [2:0] cs_tmp;
  reg [8:0] cnt;
  reg [12:0] index;               // 2^13 = 8192 > 288*18 = 5184. 18 is `data_len.  

  rom #(

  ) rom0 (
    .clk(clk),
    .addr(addr),
    .q(ramout)
  );  

  // if cs change, init = 1. not init = 0.
  always @(posedge clk) begin
    cs_tmp <= cs;
    if (cs != cs_tmp) init <= 1;
    else init <= 0;    
  end

  always @(posedge clk) begin
    if (init == 1) begin
      valid <= 0;
      index <= 0;
      cnt <= 0;
      if      (cs == `LAYER0) addr <= 0;
      else if (cs == `LAYER1) addr <= 288;
      else if (cs == `LAYER2) addr <= 2*288;
      else if (cs == `LAYER3) addr <= 3*288;
      else if (cs == `AFFINE) addr <= 4*288;
    end
    else if (cnt == 0) begin
      cnt <= cnt + 1;
      addr <= addr + 1;      
    end
    else if (cnt < 288 + 1) begin
      index <= index + `data_len;
      cnt <= cnt + 1;
      addr <= addr + 1;
    end
    else if (cnt == 288 + 1) begin
      valid <= 1;
      cnt <= cnt + 1;
    end
    q[index +: `data_len] <= ramout;
  end
  
endmodule