`include "num_data.v"

module w_rom_18 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000100011011111111111010000100000000000010011001111111111101000100000000000011010010111111111000110011111111110111100101000000000011001011111111111010001000;
    mem[1] = 162'b111111111011101111111111110111110000000000000000111011000000000010001010111111110111101000000000001100110010111111110110000010111111111101100010111111110100101001;
    mem[2] = 162'b000000000011010010111111111100010111000000000001111101111111111101111100000000000110101101111111111110100100111111111010001100111111111111110101111111111101010001;
    mem[3] = 162'b111111110101010001111111111010011101000000000010101101111111110100101000111111101111001011111111100101100000000000000010100111111111010111010000111111011110101100;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111110000011010000000001011100111111111111001111000111111111111110000000000000001000001111111111011100100111111111110001010111111111101001101111111110111001001;
    mem[33] = 162'b111111111110011110111111111101011110000000001000110100111111111100011000000000000011101001111111110101000100111111111011000111000000000111000000111111111010001101;
    mem[34] = 162'b111111110000000011111111111111101000111111111100110001111111111110010000000000000001001110000000000010000100000000000110111000111111111010011101000000000111100111;
    mem[35] = 162'b000000000000101000111111111011100001111111111100100101000000000110000100111111111101111110111111111111011001000000000010001101000000000111111101000000001000011011;
    mem[36] = 162'b000000000010001100000000000000010110111111111100000001000000000010100100000000000001110011000000001000111100000000001000111111111111111110000101000000000110101101;
    mem[37] = 162'b000000000110110010111111111001000010000000000001111011000000000001111010111111111000101101111111111111111011000000000011000010000000000010001011000000000001111101;
    mem[38] = 162'b000000000100000100000000000011101011111111111101001001000000000110010101000000000110000111000000000001001011000000001000111011000000000100001001000000001011011000;
    mem[39] = 162'b000000000101001011111111111111000100111111111011001111000000000001000001111111110111010011111111111101011110000000000101101100000000000001010001111111110110011110;
    mem[40] = 162'b000000000111111011111111111111001111000000000000100000111111111110100111000000000100010010000000001000010010000000000100110011000000000010100001111111111111010001;
    mem[41] = 162'b000000000010101000111111111001001111000000000100011101111111111010101100111111111101010011000000000010110001111111111101010110111111111011110111111111111111011011;
    mem[42] = 162'b000000000001010010111111111111101010111111111011111101111111111101101101000000000010101111000000001010101011111111111101101110111111111000111010000000001010111101;
    mem[43] = 162'b000000000001101010111111111110010000000000000001001101111111111101111110000000000000111110000000000111111000000000000100111111000000000001101011000000001001011000;
    mem[44] = 162'b111111111010001000111111111110011000111111111001000000000000000100010101111111111110110110000000000101000110000000000001111010111111111111100001111111111011000110;
    mem[45] = 162'b111111111111111011111111111110110101000000000011101000111111111110010001111111111101101101000000000000001111111111111111010101000000000001101110111111111100010111;
    mem[46] = 162'b111111111101001000111111111101000010000000000011101111111111111110111000000000001001100001111111111110001000000000000010010111111111111100111101111111111100010111;
    mem[47] = 162'b111111111011111110000000000000100111000000000011000100111111111010110110000000000110101011111111111111011001111111111010111111111111111011010011111111111100010100;
    mem[48] = 162'b111111110111010110000000000010100100000000000000110111000000000001101110000000000001101110000000000000000100000000000110001000000000000010000001111111111110111101;
    mem[49] = 162'b000000001000100010111111110011001000000000000000100010111111101110100000111111111101100011000000000010001100111111111111110000000000000000111111111111111010111100;
    mem[50] = 162'b111111111110000010111111111110011100000000000100100001111111111111110010000000000011000101000000001001100110111111111101100110111111111010010111111111111011010001;
    mem[51] = 162'b000000000111111000000000000110011100000000000110100010000000001000000000000000000110100100000000001010101000000000001000010100000000000101000010000000001010000110;
    mem[52] = 162'b000000000110001111111111111101110010000000000010110110000000000101110011000000000010101011000000000100010100000000000101011101111111111110000110000000000010110101;
    mem[53] = 162'b111111111110001101000000000101011100000000000100001101111111111111000110111111111110111111111111110111111011111111111100000111111111111111011000000000000011010011;
    mem[54] = 162'b111111111001111010000000000111111011111111111100110001000000000001010100111111111010000011111111111011101100000000000010010111111111111110011101000000000011010111;
    mem[55] = 162'b111111111111001110111111111001111100111111111110101101000000000101111111000000000010010011111111111000111001111111111101100000111111111110101100000000000000111100;
    mem[56] = 162'b000000000000101100000000000001000001111111111100101111000000001000011100111111111101101000111111111000110100000000000101100101111111111001110010111111111111110000;
    mem[57] = 162'b000000000001100101000000000001101011000000000000011000111111111110110101000000000010011111000000000001011011111111111110111111000000000001111010111111110111000000;
    mem[58] = 162'b111111111111111100111111111110110011111111111101000111000000000101110101111111111100000100000000000010000101000000000010111100000000000101011000000000000101000100;
    mem[59] = 162'b111111111100001010111111111111101000000000000111110100000000001000010001111111111100010110111111110101101100000000000010111011000000000011100101111111111111011101;
    mem[60] = 162'b111111111000110000111111110100000111000000000111110100111111111001001110111111111010110100000000000011110001111111110111101100111111111100110110000000000011110000;
    mem[61] = 162'b111111111110001111111111111110010001111111111101100011111111111010001101111111111011000101000000000001011010111111111011010110000000000000011011111111111100000011;
    mem[62] = 162'b111111111000011111111111110111111100000000000100000110000000000001110110000000000011111011111111111111010010111111111001001111111111111111100111000000000001110100;
    mem[63] = 162'b000000000100010101000000000011011111111111111110101110000000000010000001000000000010011001000000000000111111000000000000101110000000000100100010000000000000000010;
    mem[64] = 162'b000000000011111001111111111010011101000000000010011001111111111000000011000000000011111100111111111111001000000000000010100111000000000000110100111111111010100100;
    mem[65] = 162'b000000000000011110000000000000011101111111111101010110111111111101000101111111111100110010111111111011111111000000000001110110111111111111101111000000000000000100;
    mem[66] = 162'b111111111110010000111111111100100000111111111010010001000000000111110001111111111110010100111111110101010111000000001000100011111111110111100100000000000010010000;
    mem[67] = 162'b111111111111011001000000000100001110111111111011000110000000000001011000111111111101101101111111111010001001000000000100010110000000000011011000000000000001111000;
    mem[68] = 162'b000000000010001100111111111110000101111111111100001110111111111100001010000000000000111100111111111111001111111111111010100111111111111011011011111111110100010001;
    mem[69] = 162'b111111111110111100111111111101110001000000000001100000000000000011000001111111111111010101111111111100011100111111111011111001000000000100101010000000000110000000;
    mem[70] = 162'b000000000000110001111111111111110101000000000111010110111111111011101101111111111100001001000000000000111000111111111000111111000000000000011000000000000001110001;
    mem[71] = 162'b111111111100111101111111111100000110000000000001010100111111111101010010000000000000001010111111111101001011000000000101011001000000000100101011000000000101100001;
    mem[72] = 162'b000000000001101100000000000010001010000000000001101000000000000000010011111111111111010111111111111110110001111111111111001110111111111101110110000000000000001101;
    mem[73] = 162'b111111110111010001111111111101000111000000000000100111000000000001001011111111110111101100000000000010011001000000000000110010000000000000101000111111111111000100;
    mem[74] = 162'b111111111111010010111111111011011100000000000010000000111111111110110110111111111011000101000000000000001000000000000110010101111111111010111100000000000001011010;
    mem[75] = 162'b111111111111110011000000000010101001000000000001011011000000000100110011111111111110001111000000000010100001000000000110110011000000000000010101111111111010000000;
    mem[76] = 162'b000000000001000000000000000101100010111111111110100011000000000011100101000000000001100010000000000000001101000000000101110001000000001100000101000000001000010101;
    mem[77] = 162'b000000000000001101111111111110000001111111111011011001000000000000010111000000000001000101111111111101001110111111111110010101111111111011110010000000001000000010;
    mem[78] = 162'b000000000001011010000000000010111001000000000100011100000000000011110111000000001010110010000000000011110110000000000100010010000000000110011010000000000110011000;
    mem[79] = 162'b111111110111010010111111111001101000111111111101111000111111111110100001000000000101100110000000000011010111111111111010101110000000000010010101111111111100111000;
    mem[80] = 162'b000000000000101011000000000001100110111111111101111010000000000000000001000000000101010100111111111100100101000000000011110111000000000000000101000000000000001100;
    mem[81] = 162'b000000000011000001000000000000100110000000000011100001111111111111111111111111111100111000111111111110100001111111111111010111000000000001010011111111111111111010;
    mem[82] = 162'b000000000100010000111111111010011001111111111111001011000000000011010000111111111111101110111111111111100110111111111100111111000000000100010110111111111011010110;
    mem[83] = 162'b111111111111011110000000000010100001000000000010001111111111111111001010000000000001100000000000000101001001000000000000000100111111111110101011000000000101100110;
    mem[84] = 162'b000000000000000111000000000001011101111111111110000000000000000100111100000000000000001100111111111111000011111111111011100111111111111100101000111111111111001011;
    mem[85] = 162'b111111111100010010111111111100010100000000000000111100111111111011011010000000000010010001111111111111101100000000001010111101000000000101101101111111111111001110;
    mem[86] = 162'b000000000011011010111111111010010101111111111110011010000000000101000101000000000001100110000000000011001000000000000111110101000000010010110011000000001110110110;
    mem[87] = 162'b000000000010001001000000000001110011111111111011000010000000000010000000111111111101100110000000000001010000000000000000100100111111111110101010000000000011011010;
    mem[88] = 162'b000000000010011010111111111110011001000000000000111100000000000000000010000000000001110111111111111011000100111111111110011100111111111101100010111111111110101101;
    mem[89] = 162'b000000000000010100000000000001100110000000000010011011111111111111011111000000000000010111000000000100010110111111111110100011111111111010101101111111111100101101;
    mem[90] = 162'b000000000010111100000000000010000001111111111110111111000000000100011011000000000000001000111111111101011001111111111110101111111111111111110010000000000000101001;
    mem[91] = 162'b000000000000110111111111111011010001111111111110101101000000000101010111111111111101001100000000001000000001000000000110000101000000000110010101000000001001100000;
    mem[92] = 162'b111111111111001000000000000010110111000000000001011001111111111101010100000000000010100001111111110110101011111111111011110110000000000101100000000000000000100011;
    mem[93] = 162'b111111111110111010000000000000001011000000000011110111000000000011010101111111111011101000000000000001010100000000000001101001111111111110111010111111111101101001;
    mem[94] = 162'b111111111111011011111111111101100001111111111110111100111111111110100100111111111001001100000000000010011000111111111100111111111111111110110110000000000101000100;
    mem[95] = 162'b111111111100011111000000000010101111111111110111100111111111111111011000000000000010101100000000000000100111000000001000000110000000000010110110000000000001000010;
    mem[96] = 162'b000000000000001001000000000000001000000000000000000100000000000000001010000000000000001000000000000000011100000000000000000000000000000000000011000000000000010111;
    mem[97] = 162'b111111111111110111111111111111110111000000000000001011000000000000010110000000000000010110111111111111110101111111111111110101111111111111111100000000000000001010;
    mem[98] = 162'b111111111111111000111111111111110000000000000000001101000000000000010111000000000000010010111111111111110101111111111111110111111111111111101100000000000000000001;
    mem[99] = 162'b111111111111111100000000000000011100000000000000000101111111111111110100111111111111110011000000000000001011111111111111100010111111111111101101111111111111101010;
    mem[100] = 162'b000000000000001101000000000000001101000000000000011001111111111111111111111111111111111100000000000000001011000000000000001111111111111111111101000000000000000000;
    mem[101] = 162'b000000000000011110000000000000000111000000000000100011000000000000000000111111111111111010111111111111110100111111111111110110000000000000000100111111111111111110;
    mem[102] = 162'b111111111111110001000000000000000011111111111111110011111111111111111101111111111111110101111111111111111010000000000000000010000000000000000000111111111111111000;
    mem[103] = 162'b111111111111111000000000000000000001111111111111111111111111111111111101111111111111111101111111111111111011111111111111110110000000000000001100111111111111110111;
    mem[104] = 162'b000000000000011010000000000000010110111111111111110110000000000000100000000000000000001111000000000000011000000000000000001000111111111111111010000000000000001101;
    mem[105] = 162'b111111111111110001111111111111110101000000000000000100000000000000000001111111111111110011111111111111111101000000000000010111000000000000001001111111111111110001;
    mem[106] = 162'b000000000000001000000000000000010000000000000000010110000000000000001101000000000000000111000000000000010011111111111111111101000000000000000010000000000000010101;
    mem[107] = 162'b111111111111100001111111111111101101111111111111110100000000000000000011000000000000000011111111111111110001000000000000000111000000000000010100000000000000001001;
    mem[108] = 162'b000000000000000100000000000000100001000000000000001010000000000000010101000000000000000110000000000000000001000000000000000100000000000000001110000000000000001000;
    mem[109] = 162'b000000000000000111000000000000000101000000000000000100000000000000000100000000000000001100000000000000000011000000000000001111000000000000001000000000000000001010;
    mem[110] = 162'b111111111111111100000000000000000001000000000000000101111111111111111100000000000000000111000000000000001000111111111111111011000000000000000001000000000000010111;
    mem[111] = 162'b111111111111111001111111111111110011000000000000010001111111111111110001000000000000000110000000000000000101111111111111101110000000000000001010000000000000000100;
    mem[112] = 162'b000000000000011001000000000000001011000000000000101111000000000000101110111111111111111001000000000000001011000000000000000111111111111111110001000000000000011010;
    mem[113] = 162'b000000000000001000111111111111101010000000000000001010000000000000000001000000000000001111000000000000000111000000000000010000111111111111111111000000000000001111;
    mem[114] = 162'b000000000000000000000000000000000100000000000000000001111111111111111100000000000000000010000000000000000110111111111111110010111111111111111110111111111111111011;
    mem[115] = 162'b111111111111001110111111111111110101000000000000001011111111111111110011000000000000000101000000000000010101000000000000000110000000000000000110000000000000001101;
    mem[116] = 162'b111111111111111000000000000000000000000000000000000001111111111111010110000000000000000110000000000000001100000000000000000010000000000000000110111111111111110100;
    mem[117] = 162'b111111111111110001000000000000000001111111111111011011000000000000001001000000000000000110000000000000000111000000000000010000111111111111111111000000000000010111;
    mem[118] = 162'b000000000000000101111111111111110010000000000000100000000000000000000111111111111111111101000000000000000011000000000000010100000000000000011101000000000000010000;
    mem[119] = 162'b000000000000001111000000000000000001000000000000001010000000000000010000000000000000000011000000000000001111000000000000000100000000000000010011111111111111111101;
    mem[120] = 162'b111111111111111100000000000000000101111111111111111011000000000000001100111111111111111111000000000000100011111111111111111110000000000000001000111111111111101110;
    mem[121] = 162'b000000000000001100000000000000011001111111111111111111000000000000000101000000000000001010000000000000010011000000000000100010000000000000100100000000000000010101;
    mem[122] = 162'b000000000000000011111111111111111100111111111111110010000000000000011000000000000000010000111111111111111011111111111111111001111111111111110111000000000000010100;
    mem[123] = 162'b000000000000000000111111111111111101000000000000010000000000000000000100000000000000001101111111111111111100000000000000000110111111111111110011111111111111100100;
    mem[124] = 162'b000000000000001001000000000000001001111111111111110100000000000000000101000000000000000001000000000000000110000000000000000110000000000000001001000000000000010101;
    mem[125] = 162'b111111111111110101111111111111110010111111111111011110111111111111110100000000000000001001111111111111111101000000000000011001000000000000001011000000000000010001;
    mem[126] = 162'b000000000000001111111111111111110011111111111111110001111111111111111010111111111111111111111111111111111010111111111111111001000000000000001101111111111111110110;
    mem[127] = 162'b000000000000100000000000000000001001000000000000001000111111111111110000111111111111110100111111111111110000111111111111110000111111111111011001111111111111111000;
    mem[128] = 162'b000000000000001011000000000010101000000000000101000111000000000101001011111111111111100111111111111111100010000000000010000100000000000000001000000000000000010010;
    mem[129] = 162'b111111111111111110111111111111111111000000000000000101000000000000000011111111111111111111000000000000000001111111111111110111111111111111100100000000000000010010;
    mem[130] = 162'b000000000000000010000000000000001000000000000000001011000000000000001111000000000000000100000000000000000100111111111111111111000000000000000110111111111111110111;
    mem[131] = 162'b111111111111111110000000000000000111111111111111111000111111111111111100000000000000000000000000000000000000111111111111111010111111111111111010000000000000000111;
    mem[132] = 162'b111111111111101011000000000000110011111111111111101111111111111111110000000000000000100011111111111111100100000000000000001001111111111111110010111111111111100000;
    mem[133] = 162'b111111111111111101111111111111111111000000000000001101000000000000000100111111111111111110111111111111111010000000000010010110111111111111100111111111111111101111;
    mem[134] = 162'b000000000011101110000000000110000010000000000010100100000000000000000001000000000000001001000000000000000000111111111111110101000000000000001001111111111111110011;
    mem[135] = 162'b111111111111100011111111111111011111111111111111111011111111111111101100000000000000001100000000000010011111000000000001101011000000000000010101000000000100101100;
    mem[136] = 162'b000000000000000110111111111111111111111111111111110010111111111111110101111111111111110110000000000000001100000000000000000100111111111111111101000000000000000001;
    mem[137] = 162'b000000000000000000111111111111111111000000000000001010000000000000000110111111111111110111000000000000000011000000000000001000000000000000001101000000000000000001;
    mem[138] = 162'b000000000000000000000000000000000000000000000000000011000000000000001001000000000000001111000000000000001011000000000000001011000000000000000001000000000000000000;
    mem[139] = 162'b000000000000000111111111111111111110111111111111111111000000000000000100000000000000000000000000000000000000111111111111111111111111111111111111000000000000000101;
    mem[140] = 162'b000000000000010010000000000011000010000000000010111000000000000010101010000000000000000000000000000001010100111111111111000011111111111111100010111111111110001111;
    mem[141] = 162'b111111111111111101111111111111111110000000000000000100111111111111111000111111111111111100000000000000010100000000000100111000000000000001110100000000000100100011;
    mem[142] = 162'b000000000101010011000000000101011001000000000101010001111111111111101001111111111111110001111111111111101001111111111111110001111111111111110110111111111111110111;
    mem[143] = 162'b000000000001011000111111111111100100111111111110010110000000000001010111111111111111100000111111111111101100000000000000101100111111111111111100000000000011110101;
    mem[144] = 162'b111111111111111011000000000000000100111111111111111111000000000000000001111111111111111111000000000000001010000000000000001000111111111111111011111111111111111111;
    mem[145] = 162'b000000000000000011000000000000000100000000000000001011000000000000000000111111111111111010111111111111110010000000000000000011111111111111111000111111111111110110;
    mem[146] = 162'b000000000000000000000000000000001001000000000000000011000000000000001101000000000000001100000000000000000110000000000000000111000000000000000111111111111111111101;
    mem[147] = 162'b000000000000001100000000000000000011000000000000000000111111111111111100000000000000000110000000000000000111000000000000000100111111111111111110000000000000000011;
    mem[148] = 162'b111111111111110011000000000000001001000000000000000010000000000000000110111111111111111111000000000000000111000000000000001000111111111111111101111111111111111110;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000111111111111111111001;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule