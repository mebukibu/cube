`include "num_data.v"
`include "state_layer_data.v"

module add_bias (
    input wire clk,
    input wire rst_n,
    input wire load,
    input wire [3:0] cs,
    input wire [12*32*`data_len - 1:0] d,
    output reg [12*32*`data_len - 1:0] q
  );

  // use in this module
  reg [`data_len - 1:0] bias [0:32*5 - 1]; // 1 layer uses 32 bias. 5 layers.
  reg [7:0] offset;
  integer i, j;

  always @(posedge clk) begin
    if (cs == `LAYER0) offset <= 0;
    else if (cs == `LAYER1) offset <= 32;
    else if (cs == `LAYER2) offset <= 2*32;
    else if (cs == `LAYER3) offset <= 3*32;
    else if (cs == `AFFINE) offset <= 4*32;
    else offset <= 8'hXX;
  end

  always @(posedge clk, negedge rst_n) begin
    if (!rst_n) q <= 0;
    else if (load) begin
      for (i = 0; i < 32; i = i + 1) begin
        for (j = 0; j < 12; j = j + 1) begin
          q[(12*i+j)*`data_len +: `data_len] <= d[(12*i+j)*`data_len +: `data_len] + bias[i + offset];
        end
      end
    end
  end

  initial begin
    //$readmemb("data18/bias18_data.txt", bias);
    bias[0] = 18'b111111111111100101;
    bias[1] = 18'b000000000000001001;
    bias[2] = 18'b111111111011101110;
    bias[3] = 18'b111111111011101101;
    bias[4] = 18'b111111111111011010;
    bias[5] = 18'b111111111011111000;
    bias[6] = 18'b111111111011100000;
    bias[7] = 18'b000000000010110000;
    bias[8] = 18'b111111111101101010;
    bias[9] = 18'b111111111110001011;
    bias[10] = 18'b111111111111011000;
    bias[11] = 18'b111111111111001001;
    bias[12] = 18'b111111110111000001;
    bias[13] = 18'b000000000010001110;
    bias[14] = 18'b111111111110011011;
    bias[15] = 18'b000000000010111101;
    bias[16] = 18'b000000000010100111;
    bias[17] = 18'b111111111001100001;
    bias[18] = 18'b111111111011101111;
    bias[19] = 18'b111111111011111111;
    bias[20] = 18'b000000000000101101;
    bias[21] = 18'b000000000001111011;
    bias[22] = 18'b111111111110100011;
    bias[23] = 18'b111111111000111101;
    bias[24] = 18'b000000000001001011;
    bias[25] = 18'b111111111101011000;
    bias[26] = 18'b111111111100110101;
    bias[27] = 18'b111111111010101111;
    bias[28] = 18'b111111110111111101;
    bias[29] = 18'b000000000001110101;
    bias[30] = 18'b111111110110000000;
    bias[31] = 18'b111111111010110110;
    bias[32] = 18'b111111110110111110;
    bias[33] = 18'b111111110110001001;
    bias[34] = 18'b111111110001010100;
    bias[35] = 18'b111111110111011001;
    bias[36] = 18'b111111111011000101;
    bias[37] = 18'b111111110111001010;
    bias[38] = 18'b111111111001000110;
    bias[39] = 18'b111111110101010111;
    bias[40] = 18'b111111111100101000;
    bias[41] = 18'b111111111011001011;
    bias[42] = 18'b111111111010101001;
    bias[43] = 18'b111111110101110111;
    bias[44] = 18'b111111101110100100;
    bias[45] = 18'b111111111000111000;
    bias[46] = 18'b111111101111001111;
    bias[47] = 18'b111111110110011101;
    bias[48] = 18'b111111110111001100;
    bias[49] = 18'b111111110111011001;
    bias[50] = 18'b111111110101110001;
    bias[51] = 18'b111111110100000010;
    bias[52] = 18'b111111111000010110;
    bias[53] = 18'b111111110100110011;
    bias[54] = 18'b111111110011110111;
    bias[55] = 18'b111111111010100010;
    bias[56] = 18'b111111111010001100;
    bias[57] = 18'b111111111101101011;
    bias[58] = 18'b111111110101101001;
    bias[59] = 18'b111111110101010100;
    bias[60] = 18'b111111110110110100;
    bias[61] = 18'b111111111000100100;
    bias[62] = 18'b111111111010011111;
    bias[63] = 18'b111111110110111001;
    bias[64] = 18'b111111111010001010;
    bias[65] = 18'b111111110101010110;
    bias[66] = 18'b111111110111000000;
    bias[67] = 18'b111111111001000111;
    bias[68] = 18'b111111101101110110;
    bias[69] = 18'b111111110100001110;
    bias[70] = 18'b111111110001000110;
    bias[71] = 18'b111111110110010100;
    bias[72] = 18'b111111110100010101;
    bias[73] = 18'b111111111010000011;
    bias[74] = 18'b111111111100000000;
    bias[75] = 18'b111111111010010110;
    bias[76] = 18'b111111111000111001;
    bias[77] = 18'b111111111111101100;
    bias[78] = 18'b111111110111000000;
    bias[79] = 18'b111111110110110001;
    bias[80] = 18'b111111101010101110;
    bias[81] = 18'b111111111000000001;
    bias[82] = 18'b111111111001101011;
    bias[83] = 18'b111111110101001000;
    bias[84] = 18'b111111110110000010;
    bias[85] = 18'b111111110011111100;
    bias[86] = 18'b111111111100010100;
    bias[87] = 18'b111111111001100110;
    bias[88] = 18'b111111110111011001;
    bias[89] = 18'b111111101111100010;
    bias[90] = 18'b111111111101110111;
    bias[91] = 18'b111111111011101000;
    bias[92] = 18'b111111110111010100;
    bias[93] = 18'b111111111010010011;
    bias[94] = 18'b111111110110000001;
    bias[95] = 18'b111111110111100011;
    bias[96] = 18'b111111110101000000;
    bias[97] = 18'b111111111111010101;
    bias[98] = 18'b111111111111110100;
    bias[99] = 18'b111111110001001010;
    bias[100] = 18'b111111111111101000;
    bias[101] = 18'b111111110011010110;
    bias[102] = 18'b111111110010001011;
    bias[103] = 18'b111111111111110101;
    bias[104] = 18'b111111110110000011;
    bias[105] = 18'b111111111111001011;
    bias[106] = 18'b111111111111110100;
    bias[107] = 18'b111111111111101000;
    bias[108] = 18'b111111111111110110;
    bias[109] = 18'b111111111111000010;
    bias[110] = 18'b111111111111110011;
    bias[111] = 18'b111111111111011001;
    bias[112] = 18'b111111110111100100;
    bias[113] = 18'b111111111111111001;
    bias[114] = 18'b111111111111011000;
    bias[115] = 18'b111111111001110011;
    bias[116] = 18'b111111111111011001;
    bias[117] = 18'b111111101110111100;
    bias[118] = 18'b111111111111011110;
    bias[119] = 18'b111111111111010101;
    bias[120] = 18'b111111111111100110;
    bias[121] = 18'b111111111001100111;
    bias[122] = 18'b111111111111110011;
    bias[123] = 18'b111111101110100001;
    bias[124] = 18'b111111111111101111;
    bias[125] = 18'b111111111111011011;
    bias[126] = 18'b000000000000001001;
    bias[127] = 18'b111111111111001000;
    bias[128] = 18'b111111111010110001;
    bias[129] = 18'b111111111001110100;
    bias[130] = 18'b111111111011100101;
    bias[131] = 18'b111111111010001110;
    bias[132] = 18'b111111111011000101;
    bias[133] = 18'b111111111011000100;
    bias[134] = 18'b111111111010110101;
    bias[135] = 18'b111111111010000101;
    bias[136] = 18'b111111111011010010;
    bias[137] = 18'b111111111010011101;
    bias[138] = 18'b111111111010111101;
    bias[139] = 18'b111111111011011100;
    bias[140] = 18'b000000000000000000;
    bias[141] = 18'b000000000000000000;
    bias[142] = 18'b000000000000000000;
    bias[143] = 18'b000000000000000000;
    bias[144] = 18'b000000000000000000;
    bias[145] = 18'b000000000000000000;
    bias[146] = 18'b000000000000000000;
    bias[147] = 18'b000000000000000000;
    bias[148] = 18'b000000000000000000;
    bias[149] = 18'b000000000000000000;
    bias[150] = 18'b000000000000000000;
    bias[151] = 18'b000000000000000000;
    bias[152] = 18'b000000000000000000;
    bias[153] = 18'b000000000000000000;
    bias[154] = 18'b000000000000000000;
    bias[155] = 18'b000000000000000000;
    bias[156] = 18'b000000000000000000;
    bias[157] = 18'b000000000000000000;
    bias[158] = 18'b000000000000000000;
    bias[159] = 18'b000000000000000000;
  end

endmodule