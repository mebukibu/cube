`include "../data/num_data.v"

module im2col (
    input wire clk,
    input wire rst_n,
    input wire load,
    input wire [32*5*6*`data_len - 1:0] d,
    output reg valid,
    output reg [8:0] addr,
    output reg [9*`data_len - 1:0] q
  );

  reg init;

  always @(posedge clk, negedge rst_n) begin
    if (!rst_n) begin
      init <= 0;
      valid <= 0;
      addr <= 0;
      q <= 0;
    end
    else if (load) begin
      if (init) begin
        init <= 0;
        addr <= 0;
        q <= {d[12*`data_len +: 3*`data_len], d[6*`data_len +: 3*`data_len], d[0*`data_len +: 3*`data_len]};
      end
      else if (!valid) begin
        addr <= addr + 1;
        if (addr == 0) q <= {d[42*`data_len +: 3*`data_len], d[36*`data_len +: 3*`data_len], d[30*`data_len +: 3*`data_len]};
        if (addr == 1) q <= {d[72*`data_len +: 3*`data_len], d[66*`data_len +: 3*`data_len], d[60*`data_len +: 3*`data_len]};
        if (addr == 2) q <= {d[102*`data_len +: 3*`data_len], d[96*`data_len +: 3*`data_len], d[90*`data_len +: 3*`data_len]};
        if (addr == 3) q <= {d[132*`data_len +: 3*`data_len], d[126*`data_len +: 3*`data_len], d[120*`data_len +: 3*`data_len]};       
        if (addr == 4) q <= {d[162*`data_len +: 3*`data_len], d[156*`data_len +: 3*`data_len], d[150*`data_len +: 3*`data_len]};       
        if (addr == 5) q <= {d[192*`data_len +: 3*`data_len], d[186*`data_len +: 3*`data_len], d[180*`data_len +: 3*`data_len]};       
        if (addr == 6) q <= {d[222*`data_len +: 3*`data_len], d[216*`data_len +: 3*`data_len], d[210*`data_len +: 3*`data_len]};       
        if (addr == 7) q <= {d[252*`data_len +: 3*`data_len], d[246*`data_len +: 3*`data_len], d[240*`data_len +: 3*`data_len]};       
        if (addr == 8) q <= {d[282*`data_len +: 3*`data_len], d[276*`data_len +: 3*`data_len], d[270*`data_len +: 3*`data_len]};       
        if (addr == 9) q <= {d[312*`data_len +: 3*`data_len], d[306*`data_len +: 3*`data_len], d[300*`data_len +: 3*`data_len]};       
        if (addr == 10) q <= {d[342*`data_len +: 3*`data_len], d[336*`data_len +: 3*`data_len], d[330*`data_len +: 3*`data_len]};      
        if (addr == 11) q <= {d[372*`data_len +: 3*`data_len], d[366*`data_len +: 3*`data_len], d[360*`data_len +: 3*`data_len]};      
        if (addr == 12) q <= {d[402*`data_len +: 3*`data_len], d[396*`data_len +: 3*`data_len], d[390*`data_len +: 3*`data_len]};      
        if (addr == 13) q <= {d[432*`data_len +: 3*`data_len], d[426*`data_len +: 3*`data_len], d[420*`data_len +: 3*`data_len]};      
        if (addr == 14) q <= {d[462*`data_len +: 3*`data_len], d[456*`data_len +: 3*`data_len], d[450*`data_len +: 3*`data_len]};      
        if (addr == 15) q <= {d[492*`data_len +: 3*`data_len], d[486*`data_len +: 3*`data_len], d[480*`data_len +: 3*`data_len]};      
        if (addr == 16) q <= {d[522*`data_len +: 3*`data_len], d[516*`data_len +: 3*`data_len], d[510*`data_len +: 3*`data_len]};      
        if (addr == 17) q <= {d[552*`data_len +: 3*`data_len], d[546*`data_len +: 3*`data_len], d[540*`data_len +: 3*`data_len]};      
        if (addr == 18) q <= {d[582*`data_len +: 3*`data_len], d[576*`data_len +: 3*`data_len], d[570*`data_len +: 3*`data_len]};      
        if (addr == 19) q <= {d[612*`data_len +: 3*`data_len], d[606*`data_len +: 3*`data_len], d[600*`data_len +: 3*`data_len]};      
        if (addr == 20) q <= {d[642*`data_len +: 3*`data_len], d[636*`data_len +: 3*`data_len], d[630*`data_len +: 3*`data_len]};      
        if (addr == 21) q <= {d[672*`data_len +: 3*`data_len], d[666*`data_len +: 3*`data_len], d[660*`data_len +: 3*`data_len]};      
        if (addr == 22) q <= {d[702*`data_len +: 3*`data_len], d[696*`data_len +: 3*`data_len], d[690*`data_len +: 3*`data_len]};      
        if (addr == 23) q <= {d[732*`data_len +: 3*`data_len], d[726*`data_len +: 3*`data_len], d[720*`data_len +: 3*`data_len]};      
        if (addr == 24) q <= {d[762*`data_len +: 3*`data_len], d[756*`data_len +: 3*`data_len], d[750*`data_len +: 3*`data_len]};      
        if (addr == 25) q <= {d[792*`data_len +: 3*`data_len], d[786*`data_len +: 3*`data_len], d[780*`data_len +: 3*`data_len]};      
        if (addr == 26) q <= {d[822*`data_len +: 3*`data_len], d[816*`data_len +: 3*`data_len], d[810*`data_len +: 3*`data_len]};      
        if (addr == 27) q <= {d[852*`data_len +: 3*`data_len], d[846*`data_len +: 3*`data_len], d[840*`data_len +: 3*`data_len]};      
        if (addr == 28) q <= {d[882*`data_len +: 3*`data_len], d[876*`data_len +: 3*`data_len], d[870*`data_len +: 3*`data_len]};      
        if (addr == 29) q <= {d[912*`data_len +: 3*`data_len], d[906*`data_len +: 3*`data_len], d[900*`data_len +: 3*`data_len]};      
        if (addr == 30) q <= {d[942*`data_len +: 3*`data_len], d[936*`data_len +: 3*`data_len], d[930*`data_len +: 3*`data_len]};      
        if (addr == 31) q <= {d[13*`data_len +: 3*`data_len], d[7*`data_len +: 3*`data_len], d[1*`data_len +: 3*`data_len]};
        if (addr == 32) q <= {d[43*`data_len +: 3*`data_len], d[37*`data_len +: 3*`data_len], d[31*`data_len +: 3*`data_len]};
        if (addr == 33) q <= {d[73*`data_len +: 3*`data_len], d[67*`data_len +: 3*`data_len], d[61*`data_len +: 3*`data_len]};
        if (addr == 34) q <= {d[103*`data_len +: 3*`data_len], d[97*`data_len +: 3*`data_len], d[91*`data_len +: 3*`data_len]};        
        if (addr == 35) q <= {d[133*`data_len +: 3*`data_len], d[127*`data_len +: 3*`data_len], d[121*`data_len +: 3*`data_len]};      
        if (addr == 36) q <= {d[163*`data_len +: 3*`data_len], d[157*`data_len +: 3*`data_len], d[151*`data_len +: 3*`data_len]};      
        if (addr == 37) q <= {d[193*`data_len +: 3*`data_len], d[187*`data_len +: 3*`data_len], d[181*`data_len +: 3*`data_len]};      
        if (addr == 38) q <= {d[223*`data_len +: 3*`data_len], d[217*`data_len +: 3*`data_len], d[211*`data_len +: 3*`data_len]};      
        if (addr == 39) q <= {d[253*`data_len +: 3*`data_len], d[247*`data_len +: 3*`data_len], d[241*`data_len +: 3*`data_len]};
        if (addr == 40) q <= {d[283*`data_len +: 3*`data_len], d[277*`data_len +: 3*`data_len], d[271*`data_len +: 3*`data_len]};      
        if (addr == 41) q <= {d[313*`data_len +: 3*`data_len], d[307*`data_len +: 3*`data_len], d[301*`data_len +: 3*`data_len]};      
        if (addr == 42) q <= {d[343*`data_len +: 3*`data_len], d[337*`data_len +: 3*`data_len], d[331*`data_len +: 3*`data_len]};      
        if (addr == 43) q <= {d[373*`data_len +: 3*`data_len], d[367*`data_len +: 3*`data_len], d[361*`data_len +: 3*`data_len]};      
        if (addr == 44) q <= {d[403*`data_len +: 3*`data_len], d[397*`data_len +: 3*`data_len], d[391*`data_len +: 3*`data_len]};      
        if (addr == 45) q <= {d[433*`data_len +: 3*`data_len], d[427*`data_len +: 3*`data_len], d[421*`data_len +: 3*`data_len]};      
        if (addr == 46) q <= {d[463*`data_len +: 3*`data_len], d[457*`data_len +: 3*`data_len], d[451*`data_len +: 3*`data_len]};      
        if (addr == 47) q <= {d[493*`data_len +: 3*`data_len], d[487*`data_len +: 3*`data_len], d[481*`data_len +: 3*`data_len]};      
        if (addr == 48) q <= {d[523*`data_len +: 3*`data_len], d[517*`data_len +: 3*`data_len], d[511*`data_len +: 3*`data_len]};      
        if (addr == 49) q <= {d[553*`data_len +: 3*`data_len], d[547*`data_len +: 3*`data_len], d[541*`data_len +: 3*`data_len]};      
        if (addr == 50) q <= {d[583*`data_len +: 3*`data_len], d[577*`data_len +: 3*`data_len], d[571*`data_len +: 3*`data_len]};      
        if (addr == 51) q <= {d[613*`data_len +: 3*`data_len], d[607*`data_len +: 3*`data_len], d[601*`data_len +: 3*`data_len]};      
        if (addr == 52) q <= {d[643*`data_len +: 3*`data_len], d[637*`data_len +: 3*`data_len], d[631*`data_len +: 3*`data_len]};      
        if (addr == 53) q <= {d[673*`data_len +: 3*`data_len], d[667*`data_len +: 3*`data_len], d[661*`data_len +: 3*`data_len]};      
        if (addr == 54) q <= {d[703*`data_len +: 3*`data_len], d[697*`data_len +: 3*`data_len], d[691*`data_len +: 3*`data_len]};      
        if (addr == 55) q <= {d[733*`data_len +: 3*`data_len], d[727*`data_len +: 3*`data_len], d[721*`data_len +: 3*`data_len]};      
        if (addr == 56) q <= {d[763*`data_len +: 3*`data_len], d[757*`data_len +: 3*`data_len], d[751*`data_len +: 3*`data_len]};      
        if (addr == 57) q <= {d[793*`data_len +: 3*`data_len], d[787*`data_len +: 3*`data_len], d[781*`data_len +: 3*`data_len]};      
        if (addr == 58) q <= {d[823*`data_len +: 3*`data_len], d[817*`data_len +: 3*`data_len], d[811*`data_len +: 3*`data_len]};      
        if (addr == 59) q <= {d[853*`data_len +: 3*`data_len], d[847*`data_len +: 3*`data_len], d[841*`data_len +: 3*`data_len]};      
        if (addr == 60) q <= {d[883*`data_len +: 3*`data_len], d[877*`data_len +: 3*`data_len], d[871*`data_len +: 3*`data_len]};      
        if (addr == 61) q <= {d[913*`data_len +: 3*`data_len], d[907*`data_len +: 3*`data_len], d[901*`data_len +: 3*`data_len]};      
        if (addr == 62) q <= {d[943*`data_len +: 3*`data_len], d[937*`data_len +: 3*`data_len], d[931*`data_len +: 3*`data_len]};      
        if (addr == 63) q <= {d[14*`data_len +: 3*`data_len], d[8*`data_len +: 3*`data_len], d[2*`data_len +: 3*`data_len]};
        if (addr == 64) q <= {d[44*`data_len +: 3*`data_len], d[38*`data_len +: 3*`data_len], d[32*`data_len +: 3*`data_len]};
        if (addr == 65) q <= {d[74*`data_len +: 3*`data_len], d[68*`data_len +: 3*`data_len], d[62*`data_len +: 3*`data_len]};
        if (addr == 66) q <= {d[104*`data_len +: 3*`data_len], d[98*`data_len +: 3*`data_len], d[92*`data_len +: 3*`data_len]};        
        if (addr == 67) q <= {d[134*`data_len +: 3*`data_len], d[128*`data_len +: 3*`data_len], d[122*`data_len +: 3*`data_len]};      
        if (addr == 68) q <= {d[164*`data_len +: 3*`data_len], d[158*`data_len +: 3*`data_len], d[152*`data_len +: 3*`data_len]};      
        if (addr == 69) q <= {d[194*`data_len +: 3*`data_len], d[188*`data_len +: 3*`data_len], d[182*`data_len +: 3*`data_len]};      
        if (addr == 70) q <= {d[224*`data_len +: 3*`data_len], d[218*`data_len +: 3*`data_len], d[212*`data_len +: 3*`data_len]};      
        if (addr == 71) q <= {d[254*`data_len +: 3*`data_len], d[248*`data_len +: 3*`data_len], d[242*`data_len +: 3*`data_len]};      
        if (addr == 72) q <= {d[284*`data_len +: 3*`data_len], d[278*`data_len +: 3*`data_len], d[272*`data_len +: 3*`data_len]};      
        if (addr == 73) q <= {d[314*`data_len +: 3*`data_len], d[308*`data_len +: 3*`data_len], d[302*`data_len +: 3*`data_len]};      
        if (addr == 74) q <= {d[344*`data_len +: 3*`data_len], d[338*`data_len +: 3*`data_len], d[332*`data_len +: 3*`data_len]};      
        if (addr == 75) q <= {d[374*`data_len +: 3*`data_len], d[368*`data_len +: 3*`data_len], d[362*`data_len +: 3*`data_len]};      
        if (addr == 76) q <= {d[404*`data_len +: 3*`data_len], d[398*`data_len +: 3*`data_len], d[392*`data_len +: 3*`data_len]};      
        if (addr == 77) q <= {d[434*`data_len +: 3*`data_len], d[428*`data_len +: 3*`data_len], d[422*`data_len +: 3*`data_len]};      
        if (addr == 78) q <= {d[464*`data_len +: 3*`data_len], d[458*`data_len +: 3*`data_len], d[452*`data_len +: 3*`data_len]};      
        if (addr == 79) q <= {d[494*`data_len +: 3*`data_len], d[488*`data_len +: 3*`data_len], d[482*`data_len +: 3*`data_len]};      
        if (addr == 80) q <= {d[524*`data_len +: 3*`data_len], d[518*`data_len +: 3*`data_len], d[512*`data_len +: 3*`data_len]};      
        if (addr == 81) q <= {d[554*`data_len +: 3*`data_len], d[548*`data_len +: 3*`data_len], d[542*`data_len +: 3*`data_len]};      
        if (addr == 82) q <= {d[584*`data_len +: 3*`data_len], d[578*`data_len +: 3*`data_len], d[572*`data_len +: 3*`data_len]};      
        if (addr == 83) q <= {d[614*`data_len +: 3*`data_len], d[608*`data_len +: 3*`data_len], d[602*`data_len +: 3*`data_len]};      
        if (addr == 84) q <= {d[644*`data_len +: 3*`data_len], d[638*`data_len +: 3*`data_len], d[632*`data_len +: 3*`data_len]};      
        if (addr == 85) q <= {d[674*`data_len +: 3*`data_len], d[668*`data_len +: 3*`data_len], d[662*`data_len +: 3*`data_len]};      
        if (addr == 86) q <= {d[704*`data_len +: 3*`data_len], d[698*`data_len +: 3*`data_len], d[692*`data_len +: 3*`data_len]};      
        if (addr == 87) q <= {d[734*`data_len +: 3*`data_len], d[728*`data_len +: 3*`data_len], d[722*`data_len +: 3*`data_len]};      
        if (addr == 88) q <= {d[764*`data_len +: 3*`data_len], d[758*`data_len +: 3*`data_len], d[752*`data_len +: 3*`data_len]};      
        if (addr == 89) q <= {d[794*`data_len +: 3*`data_len], d[788*`data_len +: 3*`data_len], d[782*`data_len +: 3*`data_len]};      
        if (addr == 90) q <= {d[824*`data_len +: 3*`data_len], d[818*`data_len +: 3*`data_len], d[812*`data_len +: 3*`data_len]};      
        if (addr == 91) q <= {d[854*`data_len +: 3*`data_len], d[848*`data_len +: 3*`data_len], d[842*`data_len +: 3*`data_len]};      
        if (addr == 92) q <= {d[884*`data_len +: 3*`data_len], d[878*`data_len +: 3*`data_len], d[872*`data_len +: 3*`data_len]};      
        if (addr == 93) q <= {d[914*`data_len +: 3*`data_len], d[908*`data_len +: 3*`data_len], d[902*`data_len +: 3*`data_len]};      
        if (addr == 94) q <= {d[944*`data_len +: 3*`data_len], d[938*`data_len +: 3*`data_len], d[932*`data_len +: 3*`data_len]};      
        if (addr == 95) q <= {d[15*`data_len +: 3*`data_len], d[9*`data_len +: 3*`data_len], d[3*`data_len +: 3*`data_len]};
        if (addr == 96) q <= {d[45*`data_len +: 3*`data_len], d[39*`data_len +: 3*`data_len], d[33*`data_len +: 3*`data_len]};
        if (addr == 97) q <= {d[75*`data_len +: 3*`data_len], d[69*`data_len +: 3*`data_len], d[63*`data_len +: 3*`data_len]};
        if (addr == 98) q <= {d[105*`data_len +: 3*`data_len], d[99*`data_len +: 3*`data_len], d[93*`data_len +: 3*`data_len]};        
        if (addr == 99) q <= {d[135*`data_len +: 3*`data_len], d[129*`data_len +: 3*`data_len], d[123*`data_len +: 3*`data_len]};      
        if (addr == 100) q <= {d[165*`data_len +: 3*`data_len], d[159*`data_len +: 3*`data_len], d[153*`data_len +: 3*`data_len]};     
        if (addr == 101) q <= {d[195*`data_len +: 3*`data_len], d[189*`data_len +: 3*`data_len], d[183*`data_len +: 3*`data_len]};     
        if (addr == 102) q <= {d[225*`data_len +: 3*`data_len], d[219*`data_len +: 3*`data_len], d[213*`data_len +: 3*`data_len]};     
        if (addr == 103) q <= {d[255*`data_len +: 3*`data_len], d[249*`data_len +: 3*`data_len], d[243*`data_len +: 3*`data_len]};     
        if (addr == 104) q <= {d[285*`data_len +: 3*`data_len], d[279*`data_len +: 3*`data_len], d[273*`data_len +: 3*`data_len]};     
        if (addr == 105) q <= {d[315*`data_len +: 3*`data_len], d[309*`data_len +: 3*`data_len], d[303*`data_len +: 3*`data_len]};     
        if (addr == 106) q <= {d[345*`data_len +: 3*`data_len], d[339*`data_len +: 3*`data_len], d[333*`data_len +: 3*`data_len]};     
        if (addr == 107) q <= {d[375*`data_len +: 3*`data_len], d[369*`data_len +: 3*`data_len], d[363*`data_len +: 3*`data_len]};     
        if (addr == 108) q <= {d[405*`data_len +: 3*`data_len], d[399*`data_len +: 3*`data_len], d[393*`data_len +: 3*`data_len]};     
        if (addr == 109) q <= {d[435*`data_len +: 3*`data_len], d[429*`data_len +: 3*`data_len], d[423*`data_len +: 3*`data_len]};     
        if (addr == 110) q <= {d[465*`data_len +: 3*`data_len], d[459*`data_len +: 3*`data_len], d[453*`data_len +: 3*`data_len]};     
        if (addr == 111) q <= {d[495*`data_len +: 3*`data_len], d[489*`data_len +: 3*`data_len], d[483*`data_len +: 3*`data_len]};     
        if (addr == 112) q <= {d[525*`data_len +: 3*`data_len], d[519*`data_len +: 3*`data_len], d[513*`data_len +: 3*`data_len]};     
        if (addr == 113) q <= {d[555*`data_len +: 3*`data_len], d[549*`data_len +: 3*`data_len], d[543*`data_len +: 3*`data_len]};     
        if (addr == 114) q <= {d[585*`data_len +: 3*`data_len], d[579*`data_len +: 3*`data_len], d[573*`data_len +: 3*`data_len]};     
        if (addr == 115) q <= {d[615*`data_len +: 3*`data_len], d[609*`data_len +: 3*`data_len], d[603*`data_len +: 3*`data_len]};     
        if (addr == 116) q <= {d[645*`data_len +: 3*`data_len], d[639*`data_len +: 3*`data_len], d[633*`data_len +: 3*`data_len]};     
        if (addr == 117) q <= {d[675*`data_len +: 3*`data_len], d[669*`data_len +: 3*`data_len], d[663*`data_len +: 3*`data_len]};     
        if (addr == 118) q <= {d[705*`data_len +: 3*`data_len], d[699*`data_len +: 3*`data_len], d[693*`data_len +: 3*`data_len]};     
        if (addr == 119) q <= {d[735*`data_len +: 3*`data_len], d[729*`data_len +: 3*`data_len], d[723*`data_len +: 3*`data_len]};     
        if (addr == 120) q <= {d[765*`data_len +: 3*`data_len], d[759*`data_len +: 3*`data_len], d[753*`data_len +: 3*`data_len]};     
        if (addr == 121) q <= {d[795*`data_len +: 3*`data_len], d[789*`data_len +: 3*`data_len], d[783*`data_len +: 3*`data_len]};     
        if (addr == 122) q <= {d[825*`data_len +: 3*`data_len], d[819*`data_len +: 3*`data_len], d[813*`data_len +: 3*`data_len]};     
        if (addr == 123) q <= {d[855*`data_len +: 3*`data_len], d[849*`data_len +: 3*`data_len], d[843*`data_len +: 3*`data_len]};     
        if (addr == 124) q <= {d[885*`data_len +: 3*`data_len], d[879*`data_len +: 3*`data_len], d[873*`data_len +: 3*`data_len]};     
        if (addr == 125) q <= {d[915*`data_len +: 3*`data_len], d[909*`data_len +: 3*`data_len], d[903*`data_len +: 3*`data_len]};     
        if (addr == 126) q <= {d[945*`data_len +: 3*`data_len], d[939*`data_len +: 3*`data_len], d[933*`data_len +: 3*`data_len]};     
        if (addr == 127) q <= {d[18*`data_len +: 3*`data_len], d[12*`data_len +: 3*`data_len], d[6*`data_len +: 3*`data_len]};
        if (addr == 128) q <= {d[48*`data_len +: 3*`data_len], d[42*`data_len +: 3*`data_len], d[36*`data_len +: 3*`data_len]};        
        if (addr == 129) q <= {d[78*`data_len +: 3*`data_len], d[72*`data_len +: 3*`data_len], d[66*`data_len +: 3*`data_len]};        
        if (addr == 130) q <= {d[108*`data_len +: 3*`data_len], d[102*`data_len +: 3*`data_len], d[96*`data_len +: 3*`data_len]};      
        if (addr == 131) q <= {d[138*`data_len +: 3*`data_len], d[132*`data_len +: 3*`data_len], d[126*`data_len +: 3*`data_len]};     
        if (addr == 132) q <= {d[168*`data_len +: 3*`data_len], d[162*`data_len +: 3*`data_len], d[156*`data_len +: 3*`data_len]};     
        if (addr == 133) q <= {d[198*`data_len +: 3*`data_len], d[192*`data_len +: 3*`data_len], d[186*`data_len +: 3*`data_len]};     
        if (addr == 134) q <= {d[228*`data_len +: 3*`data_len], d[222*`data_len +: 3*`data_len], d[216*`data_len +: 3*`data_len]};     
        if (addr == 135) q <= {d[258*`data_len +: 3*`data_len], d[252*`data_len +: 3*`data_len], d[246*`data_len +: 3*`data_len]};     
        if (addr == 136) q <= {d[288*`data_len +: 3*`data_len], d[282*`data_len +: 3*`data_len], d[276*`data_len +: 3*`data_len]};     
        if (addr == 137) q <= {d[318*`data_len +: 3*`data_len], d[312*`data_len +: 3*`data_len], d[306*`data_len +: 3*`data_len]};     
        if (addr == 138) q <= {d[348*`data_len +: 3*`data_len], d[342*`data_len +: 3*`data_len], d[336*`data_len +: 3*`data_len]};     
        if (addr == 139) q <= {d[378*`data_len +: 3*`data_len], d[372*`data_len +: 3*`data_len], d[366*`data_len +: 3*`data_len]};     
        if (addr == 140) q <= {d[408*`data_len +: 3*`data_len], d[402*`data_len +: 3*`data_len], d[396*`data_len +: 3*`data_len]};     
        if (addr == 141) q <= {d[438*`data_len +: 3*`data_len], d[432*`data_len +: 3*`data_len], d[426*`data_len +: 3*`data_len]};     
        if (addr == 142) q <= {d[468*`data_len +: 3*`data_len], d[462*`data_len +: 3*`data_len], d[456*`data_len +: 3*`data_len]};     
        if (addr == 143) q <= {d[498*`data_len +: 3*`data_len], d[492*`data_len +: 3*`data_len], d[486*`data_len +: 3*`data_len]};     
        if (addr == 144) q <= {d[528*`data_len +: 3*`data_len], d[522*`data_len +: 3*`data_len], d[516*`data_len +: 3*`data_len]};     
        if (addr == 145) q <= {d[558*`data_len +: 3*`data_len], d[552*`data_len +: 3*`data_len], d[546*`data_len +: 3*`data_len]};     
        if (addr == 146) q <= {d[588*`data_len +: 3*`data_len], d[582*`data_len +: 3*`data_len], d[576*`data_len +: 3*`data_len]};     
        if (addr == 147) q <= {d[618*`data_len +: 3*`data_len], d[612*`data_len +: 3*`data_len], d[606*`data_len +: 3*`data_len]};     
        if (addr == 148) q <= {d[648*`data_len +: 3*`data_len], d[642*`data_len +: 3*`data_len], d[636*`data_len +: 3*`data_len]};     
        if (addr == 149) q <= {d[678*`data_len +: 3*`data_len], d[672*`data_len +: 3*`data_len], d[666*`data_len +: 3*`data_len]};     
        if (addr == 150) q <= {d[708*`data_len +: 3*`data_len], d[702*`data_len +: 3*`data_len], d[696*`data_len +: 3*`data_len]};     
        if (addr == 151) q <= {d[738*`data_len +: 3*`data_len], d[732*`data_len +: 3*`data_len], d[726*`data_len +: 3*`data_len]};     
        if (addr == 152) q <= {d[768*`data_len +: 3*`data_len], d[762*`data_len +: 3*`data_len], d[756*`data_len +: 3*`data_len]};     
        if (addr == 153) q <= {d[798*`data_len +: 3*`data_len], d[792*`data_len +: 3*`data_len], d[786*`data_len +: 3*`data_len]};     
        if (addr == 154) q <= {d[828*`data_len +: 3*`data_len], d[822*`data_len +: 3*`data_len], d[816*`data_len +: 3*`data_len]};     
        if (addr == 155) q <= {d[858*`data_len +: 3*`data_len], d[852*`data_len +: 3*`data_len], d[846*`data_len +: 3*`data_len]};     
        if (addr == 156) q <= {d[888*`data_len +: 3*`data_len], d[882*`data_len +: 3*`data_len], d[876*`data_len +: 3*`data_len]};     
        if (addr == 157) q <= {d[918*`data_len +: 3*`data_len], d[912*`data_len +: 3*`data_len], d[906*`data_len +: 3*`data_len]};     
        if (addr == 158) q <= {d[948*`data_len +: 3*`data_len], d[942*`data_len +: 3*`data_len], d[936*`data_len +: 3*`data_len]};
        if (addr == 159) q <= {d[19*`data_len +: 3*`data_len], d[13*`data_len +: 3*`data_len], d[7*`data_len +: 3*`data_len]};
        if (addr == 160) q <= {d[49*`data_len +: 3*`data_len], d[43*`data_len +: 3*`data_len], d[37*`data_len +: 3*`data_len]};        
        if (addr == 161) q <= {d[79*`data_len +: 3*`data_len], d[73*`data_len +: 3*`data_len], d[67*`data_len +: 3*`data_len]};        
        if (addr == 162) q <= {d[109*`data_len +: 3*`data_len], d[103*`data_len +: 3*`data_len], d[97*`data_len +: 3*`data_len]};      
        if (addr == 163) q <= {d[139*`data_len +: 3*`data_len], d[133*`data_len +: 3*`data_len], d[127*`data_len +: 3*`data_len]};     
        if (addr == 164) q <= {d[169*`data_len +: 3*`data_len], d[163*`data_len +: 3*`data_len], d[157*`data_len +: 3*`data_len]};     
        if (addr == 165) q <= {d[199*`data_len +: 3*`data_len], d[193*`data_len +: 3*`data_len], d[187*`data_len +: 3*`data_len]};     
        if (addr == 166) q <= {d[229*`data_len +: 3*`data_len], d[223*`data_len +: 3*`data_len], d[217*`data_len +: 3*`data_len]};     
        if (addr == 167) q <= {d[259*`data_len +: 3*`data_len], d[253*`data_len +: 3*`data_len], d[247*`data_len +: 3*`data_len]};     
        if (addr == 168) q <= {d[289*`data_len +: 3*`data_len], d[283*`data_len +: 3*`data_len], d[277*`data_len +: 3*`data_len]};     
        if (addr == 169) q <= {d[319*`data_len +: 3*`data_len], d[313*`data_len +: 3*`data_len], d[307*`data_len +: 3*`data_len]};     
        if (addr == 170) q <= {d[349*`data_len +: 3*`data_len], d[343*`data_len +: 3*`data_len], d[337*`data_len +: 3*`data_len]};     
        if (addr == 171) q <= {d[379*`data_len +: 3*`data_len], d[373*`data_len +: 3*`data_len], d[367*`data_len +: 3*`data_len]};     
        if (addr == 172) q <= {d[409*`data_len +: 3*`data_len], d[403*`data_len +: 3*`data_len], d[397*`data_len +: 3*`data_len]};     
        if (addr == 173) q <= {d[439*`data_len +: 3*`data_len], d[433*`data_len +: 3*`data_len], d[427*`data_len +: 3*`data_len]};     
        if (addr == 174) q <= {d[469*`data_len +: 3*`data_len], d[463*`data_len +: 3*`data_len], d[457*`data_len +: 3*`data_len]};     
        if (addr == 175) q <= {d[499*`data_len +: 3*`data_len], d[493*`data_len +: 3*`data_len], d[487*`data_len +: 3*`data_len]};     
        if (addr == 176) q <= {d[529*`data_len +: 3*`data_len], d[523*`data_len +: 3*`data_len], d[517*`data_len +: 3*`data_len]};     
        if (addr == 177) q <= {d[559*`data_len +: 3*`data_len], d[553*`data_len +: 3*`data_len], d[547*`data_len +: 3*`data_len]};     
        if (addr == 178) q <= {d[589*`data_len +: 3*`data_len], d[583*`data_len +: 3*`data_len], d[577*`data_len +: 3*`data_len]};     
        if (addr == 179) q <= {d[619*`data_len +: 3*`data_len], d[613*`data_len +: 3*`data_len], d[607*`data_len +: 3*`data_len]};     
        if (addr == 180) q <= {d[649*`data_len +: 3*`data_len], d[643*`data_len +: 3*`data_len], d[637*`data_len +: 3*`data_len]};     
        if (addr == 181) q <= {d[679*`data_len +: 3*`data_len], d[673*`data_len +: 3*`data_len], d[667*`data_len +: 3*`data_len]};     
        if (addr == 182) q <= {d[709*`data_len +: 3*`data_len], d[703*`data_len +: 3*`data_len], d[697*`data_len +: 3*`data_len]};     
        if (addr == 183) q <= {d[739*`data_len +: 3*`data_len], d[733*`data_len +: 3*`data_len], d[727*`data_len +: 3*`data_len]};     
        if (addr == 184) q <= {d[769*`data_len +: 3*`data_len], d[763*`data_len +: 3*`data_len], d[757*`data_len +: 3*`data_len]};     
        if (addr == 185) q <= {d[799*`data_len +: 3*`data_len], d[793*`data_len +: 3*`data_len], d[787*`data_len +: 3*`data_len]};     
        if (addr == 186) q <= {d[829*`data_len +: 3*`data_len], d[823*`data_len +: 3*`data_len], d[817*`data_len +: 3*`data_len]};     
        if (addr == 187) q <= {d[859*`data_len +: 3*`data_len], d[853*`data_len +: 3*`data_len], d[847*`data_len +: 3*`data_len]};     
        if (addr == 188) q <= {d[889*`data_len +: 3*`data_len], d[883*`data_len +: 3*`data_len], d[877*`data_len +: 3*`data_len]};     
        if (addr == 189) q <= {d[919*`data_len +: 3*`data_len], d[913*`data_len +: 3*`data_len], d[907*`data_len +: 3*`data_len]};     
        if (addr == 190) q <= {d[949*`data_len +: 3*`data_len], d[943*`data_len +: 3*`data_len], d[937*`data_len +: 3*`data_len]};     
        if (addr == 191) q <= {d[20*`data_len +: 3*`data_len], d[14*`data_len +: 3*`data_len], d[8*`data_len +: 3*`data_len]};
        if (addr == 192) q <= {d[50*`data_len +: 3*`data_len], d[44*`data_len +: 3*`data_len], d[38*`data_len +: 3*`data_len]};        
        if (addr == 193) q <= {d[80*`data_len +: 3*`data_len], d[74*`data_len +: 3*`data_len], d[68*`data_len +: 3*`data_len]};        
        if (addr == 194) q <= {d[110*`data_len +: 3*`data_len], d[104*`data_len +: 3*`data_len], d[98*`data_len +: 3*`data_len]};      
        if (addr == 195) q <= {d[140*`data_len +: 3*`data_len], d[134*`data_len +: 3*`data_len], d[128*`data_len +: 3*`data_len]};     
        if (addr == 196) q <= {d[170*`data_len +: 3*`data_len], d[164*`data_len +: 3*`data_len], d[158*`data_len +: 3*`data_len]};     
        if (addr == 197) q <= {d[200*`data_len +: 3*`data_len], d[194*`data_len +: 3*`data_len], d[188*`data_len +: 3*`data_len]};     
        if (addr == 198) q <= {d[230*`data_len +: 3*`data_len], d[224*`data_len +: 3*`data_len], d[218*`data_len +: 3*`data_len]};     
        if (addr == 199) q <= {d[260*`data_len +: 3*`data_len], d[254*`data_len +: 3*`data_len], d[248*`data_len +: 3*`data_len]};     
        if (addr == 200) q <= {d[290*`data_len +: 3*`data_len], d[284*`data_len +: 3*`data_len], d[278*`data_len +: 3*`data_len]};     
        if (addr == 201) q <= {d[320*`data_len +: 3*`data_len], d[314*`data_len +: 3*`data_len], d[308*`data_len +: 3*`data_len]};     
        if (addr == 202) q <= {d[350*`data_len +: 3*`data_len], d[344*`data_len +: 3*`data_len], d[338*`data_len +: 3*`data_len]};     
        if (addr == 203) q <= {d[380*`data_len +: 3*`data_len], d[374*`data_len +: 3*`data_len], d[368*`data_len +: 3*`data_len]};     
        if (addr == 204) q <= {d[410*`data_len +: 3*`data_len], d[404*`data_len +: 3*`data_len], d[398*`data_len +: 3*`data_len]};     
        if (addr == 205) q <= {d[440*`data_len +: 3*`data_len], d[434*`data_len +: 3*`data_len], d[428*`data_len +: 3*`data_len]};     
        if (addr == 206) q <= {d[470*`data_len +: 3*`data_len], d[464*`data_len +: 3*`data_len], d[458*`data_len +: 3*`data_len]};     
        if (addr == 207) q <= {d[500*`data_len +: 3*`data_len], d[494*`data_len +: 3*`data_len], d[488*`data_len +: 3*`data_len]};     
        if (addr == 208) q <= {d[530*`data_len +: 3*`data_len], d[524*`data_len +: 3*`data_len], d[518*`data_len +: 3*`data_len]};     
        if (addr == 209) q <= {d[560*`data_len +: 3*`data_len], d[554*`data_len +: 3*`data_len], d[548*`data_len +: 3*`data_len]};     
        if (addr == 210) q <= {d[590*`data_len +: 3*`data_len], d[584*`data_len +: 3*`data_len], d[578*`data_len +: 3*`data_len]};     
        if (addr == 211) q <= {d[620*`data_len +: 3*`data_len], d[614*`data_len +: 3*`data_len], d[608*`data_len +: 3*`data_len]};     
        if (addr == 212) q <= {d[650*`data_len +: 3*`data_len], d[644*`data_len +: 3*`data_len], d[638*`data_len +: 3*`data_len]};
        if (addr == 213) q <= {d[680*`data_len +: 3*`data_len], d[674*`data_len +: 3*`data_len], d[668*`data_len +: 3*`data_len]};     
        if (addr == 214) q <= {d[710*`data_len +: 3*`data_len], d[704*`data_len +: 3*`data_len], d[698*`data_len +: 3*`data_len]};     
        if (addr == 215) q <= {d[740*`data_len +: 3*`data_len], d[734*`data_len +: 3*`data_len], d[728*`data_len +: 3*`data_len]};     
        if (addr == 216) q <= {d[770*`data_len +: 3*`data_len], d[764*`data_len +: 3*`data_len], d[758*`data_len +: 3*`data_len]};     
        if (addr == 217) q <= {d[800*`data_len +: 3*`data_len], d[794*`data_len +: 3*`data_len], d[788*`data_len +: 3*`data_len]};     
        if (addr == 218) q <= {d[830*`data_len +: 3*`data_len], d[824*`data_len +: 3*`data_len], d[818*`data_len +: 3*`data_len]};     
        if (addr == 219) q <= {d[860*`data_len +: 3*`data_len], d[854*`data_len +: 3*`data_len], d[848*`data_len +: 3*`data_len]};     
        if (addr == 220) q <= {d[890*`data_len +: 3*`data_len], d[884*`data_len +: 3*`data_len], d[878*`data_len +: 3*`data_len]};     
        if (addr == 221) q <= {d[920*`data_len +: 3*`data_len], d[914*`data_len +: 3*`data_len], d[908*`data_len +: 3*`data_len]};     
        if (addr == 222) q <= {d[950*`data_len +: 3*`data_len], d[944*`data_len +: 3*`data_len], d[938*`data_len +: 3*`data_len]};     
        if (addr == 223) q <= {d[21*`data_len +: 3*`data_len], d[15*`data_len +: 3*`data_len], d[9*`data_len +: 3*`data_len]};
        if (addr == 224) q <= {d[51*`data_len +: 3*`data_len], d[45*`data_len +: 3*`data_len], d[39*`data_len +: 3*`data_len]};        
        if (addr == 225) q <= {d[81*`data_len +: 3*`data_len], d[75*`data_len +: 3*`data_len], d[69*`data_len +: 3*`data_len]};        
        if (addr == 226) q <= {d[111*`data_len +: 3*`data_len], d[105*`data_len +: 3*`data_len], d[99*`data_len +: 3*`data_len]};      
        if (addr == 227) q <= {d[141*`data_len +: 3*`data_len], d[135*`data_len +: 3*`data_len], d[129*`data_len +: 3*`data_len]};     
        if (addr == 228) q <= {d[171*`data_len +: 3*`data_len], d[165*`data_len +: 3*`data_len], d[159*`data_len +: 3*`data_len]};     
        if (addr == 229) q <= {d[201*`data_len +: 3*`data_len], d[195*`data_len +: 3*`data_len], d[189*`data_len +: 3*`data_len]};     
        if (addr == 230) q <= {d[231*`data_len +: 3*`data_len], d[225*`data_len +: 3*`data_len], d[219*`data_len +: 3*`data_len]};     
        if (addr == 231) q <= {d[261*`data_len +: 3*`data_len], d[255*`data_len +: 3*`data_len], d[249*`data_len +: 3*`data_len]};     
        if (addr == 232) q <= {d[291*`data_len +: 3*`data_len], d[285*`data_len +: 3*`data_len], d[279*`data_len +: 3*`data_len]};     
        if (addr == 233) q <= {d[321*`data_len +: 3*`data_len], d[315*`data_len +: 3*`data_len], d[309*`data_len +: 3*`data_len]};     
        if (addr == 234) q <= {d[351*`data_len +: 3*`data_len], d[345*`data_len +: 3*`data_len], d[339*`data_len +: 3*`data_len]};     
        if (addr == 235) q <= {d[381*`data_len +: 3*`data_len], d[375*`data_len +: 3*`data_len], d[369*`data_len +: 3*`data_len]};     
        if (addr == 236) q <= {d[411*`data_len +: 3*`data_len], d[405*`data_len +: 3*`data_len], d[399*`data_len +: 3*`data_len]};     
        if (addr == 237) q <= {d[441*`data_len +: 3*`data_len], d[435*`data_len +: 3*`data_len], d[429*`data_len +: 3*`data_len]};     
        if (addr == 238) q <= {d[471*`data_len +: 3*`data_len], d[465*`data_len +: 3*`data_len], d[459*`data_len +: 3*`data_len]};     
        if (addr == 239) q <= {d[501*`data_len +: 3*`data_len], d[495*`data_len +: 3*`data_len], d[489*`data_len +: 3*`data_len]};     
        if (addr == 240) q <= {d[531*`data_len +: 3*`data_len], d[525*`data_len +: 3*`data_len], d[519*`data_len +: 3*`data_len]};     
        if (addr == 241) q <= {d[561*`data_len +: 3*`data_len], d[555*`data_len +: 3*`data_len], d[549*`data_len +: 3*`data_len]};     
        if (addr == 242) q <= {d[591*`data_len +: 3*`data_len], d[585*`data_len +: 3*`data_len], d[579*`data_len +: 3*`data_len]};     
        if (addr == 243) q <= {d[621*`data_len +: 3*`data_len], d[615*`data_len +: 3*`data_len], d[609*`data_len +: 3*`data_len]};     
        if (addr == 244) q <= {d[651*`data_len +: 3*`data_len], d[645*`data_len +: 3*`data_len], d[639*`data_len +: 3*`data_len]};     
        if (addr == 245) q <= {d[681*`data_len +: 3*`data_len], d[675*`data_len +: 3*`data_len], d[669*`data_len +: 3*`data_len]};     
        if (addr == 246) q <= {d[711*`data_len +: 3*`data_len], d[705*`data_len +: 3*`data_len], d[699*`data_len +: 3*`data_len]};     
        if (addr == 247) q <= {d[741*`data_len +: 3*`data_len], d[735*`data_len +: 3*`data_len], d[729*`data_len +: 3*`data_len]};     
        if (addr == 248) q <= {d[771*`data_len +: 3*`data_len], d[765*`data_len +: 3*`data_len], d[759*`data_len +: 3*`data_len]};     
        if (addr == 249) q <= {d[801*`data_len +: 3*`data_len], d[795*`data_len +: 3*`data_len], d[789*`data_len +: 3*`data_len]};     
        if (addr == 250) q <= {d[831*`data_len +: 3*`data_len], d[825*`data_len +: 3*`data_len], d[819*`data_len +: 3*`data_len]};     
        if (addr == 251) q <= {d[861*`data_len +: 3*`data_len], d[855*`data_len +: 3*`data_len], d[849*`data_len +: 3*`data_len]};     
        if (addr == 252) q <= {d[891*`data_len +: 3*`data_len], d[885*`data_len +: 3*`data_len], d[879*`data_len +: 3*`data_len]};     
        if (addr == 253) q <= {d[921*`data_len +: 3*`data_len], d[915*`data_len +: 3*`data_len], d[909*`data_len +: 3*`data_len]};     
        if (addr == 254) q <= {d[951*`data_len +: 3*`data_len], d[945*`data_len +: 3*`data_len], d[939*`data_len +: 3*`data_len]};     
        if (addr == 255) q <= {d[24*`data_len +: 3*`data_len], d[18*`data_len +: 3*`data_len], d[12*`data_len +: 3*`data_len]};        
        if (addr == 256) q <= {d[54*`data_len +: 3*`data_len], d[48*`data_len +: 3*`data_len], d[42*`data_len +: 3*`data_len]};        
        if (addr == 257) q <= {d[84*`data_len +: 3*`data_len], d[78*`data_len +: 3*`data_len], d[72*`data_len +: 3*`data_len]};        
        if (addr == 258) q <= {d[114*`data_len +: 3*`data_len], d[108*`data_len +: 3*`data_len], d[102*`data_len +: 3*`data_len]};     
        if (addr == 259) q <= {d[144*`data_len +: 3*`data_len], d[138*`data_len +: 3*`data_len], d[132*`data_len +: 3*`data_len]};     
        if (addr == 260) q <= {d[174*`data_len +: 3*`data_len], d[168*`data_len +: 3*`data_len], d[162*`data_len +: 3*`data_len]};     
        if (addr == 261) q <= {d[204*`data_len +: 3*`data_len], d[198*`data_len +: 3*`data_len], d[192*`data_len +: 3*`data_len]};     
        if (addr == 262) q <= {d[234*`data_len +: 3*`data_len], d[228*`data_len +: 3*`data_len], d[222*`data_len +: 3*`data_len]};     
        if (addr == 263) q <= {d[264*`data_len +: 3*`data_len], d[258*`data_len +: 3*`data_len], d[252*`data_len +: 3*`data_len]};     
        if (addr == 264) q <= {d[294*`data_len +: 3*`data_len], d[288*`data_len +: 3*`data_len], d[282*`data_len +: 3*`data_len]};     
        if (addr == 265) q <= {d[324*`data_len +: 3*`data_len], d[318*`data_len +: 3*`data_len], d[312*`data_len +: 3*`data_len]};     
        if (addr == 266) q <= {d[354*`data_len +: 3*`data_len], d[348*`data_len +: 3*`data_len], d[342*`data_len +: 3*`data_len]};     
        if (addr == 267) q <= {d[384*`data_len +: 3*`data_len], d[378*`data_len +: 3*`data_len], d[372*`data_len +: 3*`data_len]};     
        if (addr == 268) q <= {d[414*`data_len +: 3*`data_len], d[408*`data_len +: 3*`data_len], d[402*`data_len +: 3*`data_len]};     
        if (addr == 269) q <= {d[444*`data_len +: 3*`data_len], d[438*`data_len +: 3*`data_len], d[432*`data_len +: 3*`data_len]};     
        if (addr == 270) q <= {d[474*`data_len +: 3*`data_len], d[468*`data_len +: 3*`data_len], d[462*`data_len +: 3*`data_len]};     
        if (addr == 271) q <= {d[504*`data_len +: 3*`data_len], d[498*`data_len +: 3*`data_len], d[492*`data_len +: 3*`data_len]};     
        if (addr == 272) q <= {d[534*`data_len +: 3*`data_len], d[528*`data_len +: 3*`data_len], d[522*`data_len +: 3*`data_len]};     
        if (addr == 273) q <= {d[564*`data_len +: 3*`data_len], d[558*`data_len +: 3*`data_len], d[552*`data_len +: 3*`data_len]};     
        if (addr == 274) q <= {d[594*`data_len +: 3*`data_len], d[588*`data_len +: 3*`data_len], d[582*`data_len +: 3*`data_len]};     
        if (addr == 275) q <= {d[624*`data_len +: 3*`data_len], d[618*`data_len +: 3*`data_len], d[612*`data_len +: 3*`data_len]};
        if (addr == 276) q <= {d[654*`data_len +: 3*`data_len], d[648*`data_len +: 3*`data_len], d[642*`data_len +: 3*`data_len]};     
        if (addr == 277) q <= {d[684*`data_len +: 3*`data_len], d[678*`data_len +: 3*`data_len], d[672*`data_len +: 3*`data_len]};     
        if (addr == 278) q <= {d[714*`data_len +: 3*`data_len], d[708*`data_len +: 3*`data_len], d[702*`data_len +: 3*`data_len]};     
        if (addr == 279) q <= {d[744*`data_len +: 3*`data_len], d[738*`data_len +: 3*`data_len], d[732*`data_len +: 3*`data_len]};     
        if (addr == 280) q <= {d[774*`data_len +: 3*`data_len], d[768*`data_len +: 3*`data_len], d[762*`data_len +: 3*`data_len]};     
        if (addr == 281) q <= {d[804*`data_len +: 3*`data_len], d[798*`data_len +: 3*`data_len], d[792*`data_len +: 3*`data_len]};     
        if (addr == 282) q <= {d[834*`data_len +: 3*`data_len], d[828*`data_len +: 3*`data_len], d[822*`data_len +: 3*`data_len]};     
        if (addr == 283) q <= {d[864*`data_len +: 3*`data_len], d[858*`data_len +: 3*`data_len], d[852*`data_len +: 3*`data_len]};     
        if (addr == 284) q <= {d[894*`data_len +: 3*`data_len], d[888*`data_len +: 3*`data_len], d[882*`data_len +: 3*`data_len]};     
        if (addr == 285) q <= {d[924*`data_len +: 3*`data_len], d[918*`data_len +: 3*`data_len], d[912*`data_len +: 3*`data_len]};     
        if (addr == 286) q <= {d[954*`data_len +: 3*`data_len], d[948*`data_len +: 3*`data_len], d[942*`data_len +: 3*`data_len]};     
        if (addr == 287) q <= {d[25*`data_len +: 3*`data_len], d[19*`data_len +: 3*`data_len], d[13*`data_len +: 3*`data_len]};        
        if (addr == 288) q <= {d[55*`data_len +: 3*`data_len], d[49*`data_len +: 3*`data_len], d[43*`data_len +: 3*`data_len]};        
        if (addr == 289) q <= {d[85*`data_len +: 3*`data_len], d[79*`data_len +: 3*`data_len], d[73*`data_len +: 3*`data_len]};        
        if (addr == 290) q <= {d[115*`data_len +: 3*`data_len], d[109*`data_len +: 3*`data_len], d[103*`data_len +: 3*`data_len]};     
        if (addr == 291) q <= {d[145*`data_len +: 3*`data_len], d[139*`data_len +: 3*`data_len], d[133*`data_len +: 3*`data_len]};     
        if (addr == 292) q <= {d[175*`data_len +: 3*`data_len], d[169*`data_len +: 3*`data_len], d[163*`data_len +: 3*`data_len]};     
        if (addr == 293) q <= {d[205*`data_len +: 3*`data_len], d[199*`data_len +: 3*`data_len], d[193*`data_len +: 3*`data_len]};     
        if (addr == 294) q <= {d[235*`data_len +: 3*`data_len], d[229*`data_len +: 3*`data_len], d[223*`data_len +: 3*`data_len]};     
        if (addr == 295) q <= {d[265*`data_len +: 3*`data_len], d[259*`data_len +: 3*`data_len], d[253*`data_len +: 3*`data_len]};     
        if (addr == 296) q <= {d[295*`data_len +: 3*`data_len], d[289*`data_len +: 3*`data_len], d[283*`data_len +: 3*`data_len]};     
        if (addr == 297) q <= {d[325*`data_len +: 3*`data_len], d[319*`data_len +: 3*`data_len], d[313*`data_len +: 3*`data_len]};     
        if (addr == 298) q <= {d[355*`data_len +: 3*`data_len], d[349*`data_len +: 3*`data_len], d[343*`data_len +: 3*`data_len]};     
        if (addr == 299) q <= {d[385*`data_len +: 3*`data_len], d[379*`data_len +: 3*`data_len], d[373*`data_len +: 3*`data_len]};     
        if (addr == 300) q <= {d[415*`data_len +: 3*`data_len], d[409*`data_len +: 3*`data_len], d[403*`data_len +: 3*`data_len]};     
        if (addr == 301) q <= {d[445*`data_len +: 3*`data_len], d[439*`data_len +: 3*`data_len], d[433*`data_len +: 3*`data_len]};     
        if (addr == 302) q <= {d[475*`data_len +: 3*`data_len], d[469*`data_len +: 3*`data_len], d[463*`data_len +: 3*`data_len]};     
        if (addr == 303) q <= {d[505*`data_len +: 3*`data_len], d[499*`data_len +: 3*`data_len], d[493*`data_len +: 3*`data_len]};     
        if (addr == 304) q <= {d[535*`data_len +: 3*`data_len], d[529*`data_len +: 3*`data_len], d[523*`data_len +: 3*`data_len]};     
        if (addr == 305) q <= {d[565*`data_len +: 3*`data_len], d[559*`data_len +: 3*`data_len], d[553*`data_len +: 3*`data_len]};     
        if (addr == 306) q <= {d[595*`data_len +: 3*`data_len], d[589*`data_len +: 3*`data_len], d[583*`data_len +: 3*`data_len]};     
        if (addr == 307) q <= {d[625*`data_len +: 3*`data_len], d[619*`data_len +: 3*`data_len], d[613*`data_len +: 3*`data_len]};     
        if (addr == 308) q <= {d[655*`data_len +: 3*`data_len], d[649*`data_len +: 3*`data_len], d[643*`data_len +: 3*`data_len]};     
        if (addr == 309) q <= {d[685*`data_len +: 3*`data_len], d[679*`data_len +: 3*`data_len], d[673*`data_len +: 3*`data_len]};     
        if (addr == 310) q <= {d[715*`data_len +: 3*`data_len], d[709*`data_len +: 3*`data_len], d[703*`data_len +: 3*`data_len]};     
        if (addr == 311) q <= {d[745*`data_len +: 3*`data_len], d[739*`data_len +: 3*`data_len], d[733*`data_len +: 3*`data_len]};     
        if (addr == 312) q <= {d[775*`data_len +: 3*`data_len], d[769*`data_len +: 3*`data_len], d[763*`data_len +: 3*`data_len]};     
        if (addr == 313) q <= {d[805*`data_len +: 3*`data_len], d[799*`data_len +: 3*`data_len], d[793*`data_len +: 3*`data_len]};     
        if (addr == 314) q <= {d[835*`data_len +: 3*`data_len], d[829*`data_len +: 3*`data_len], d[823*`data_len +: 3*`data_len]};     
        if (addr == 315) q <= {d[865*`data_len +: 3*`data_len], d[859*`data_len +: 3*`data_len], d[853*`data_len +: 3*`data_len]};     
        if (addr == 316) q <= {d[895*`data_len +: 3*`data_len], d[889*`data_len +: 3*`data_len], d[883*`data_len +: 3*`data_len]};     
        if (addr == 317) q <= {d[925*`data_len +: 3*`data_len], d[919*`data_len +: 3*`data_len], d[913*`data_len +: 3*`data_len]};     
        if (addr == 318) q <= {d[955*`data_len +: 3*`data_len], d[949*`data_len +: 3*`data_len], d[943*`data_len +: 3*`data_len]};     
        if (addr == 319) q <= {d[26*`data_len +: 3*`data_len], d[20*`data_len +: 3*`data_len], d[14*`data_len +: 3*`data_len]};        
        if (addr == 320) q <= {d[56*`data_len +: 3*`data_len], d[50*`data_len +: 3*`data_len], d[44*`data_len +: 3*`data_len]};        
        if (addr == 321) q <= {d[86*`data_len +: 3*`data_len], d[80*`data_len +: 3*`data_len], d[74*`data_len +: 3*`data_len]};        
        if (addr == 322) q <= {d[116*`data_len +: 3*`data_len], d[110*`data_len +: 3*`data_len], d[104*`data_len +: 3*`data_len]};     
        if (addr == 323) q <= {d[146*`data_len +: 3*`data_len], d[140*`data_len +: 3*`data_len], d[134*`data_len +: 3*`data_len]};     
        if (addr == 324) q <= {d[176*`data_len +: 3*`data_len], d[170*`data_len +: 3*`data_len], d[164*`data_len +: 3*`data_len]};     
        if (addr == 325) q <= {d[206*`data_len +: 3*`data_len], d[200*`data_len +: 3*`data_len], d[194*`data_len +: 3*`data_len]};     
        if (addr == 326) q <= {d[236*`data_len +: 3*`data_len], d[230*`data_len +: 3*`data_len], d[224*`data_len +: 3*`data_len]};     
        if (addr == 327) q <= {d[266*`data_len +: 3*`data_len], d[260*`data_len +: 3*`data_len], d[254*`data_len +: 3*`data_len]};     
        if (addr == 328) q <= {d[296*`data_len +: 3*`data_len], d[290*`data_len +: 3*`data_len], d[284*`data_len +: 3*`data_len]};     
        if (addr == 329) q <= {d[326*`data_len +: 3*`data_len], d[320*`data_len +: 3*`data_len], d[314*`data_len +: 3*`data_len]};     
        if (addr == 330) q <= {d[356*`data_len +: 3*`data_len], d[350*`data_len +: 3*`data_len], d[344*`data_len +: 3*`data_len]};     
        if (addr == 331) q <= {d[386*`data_len +: 3*`data_len], d[380*`data_len +: 3*`data_len], d[374*`data_len +: 3*`data_len]};     
        if (addr == 332) q <= {d[416*`data_len +: 3*`data_len], d[410*`data_len +: 3*`data_len], d[404*`data_len +: 3*`data_len]};     
        if (addr == 333) q <= {d[446*`data_len +: 3*`data_len], d[440*`data_len +: 3*`data_len], d[434*`data_len +: 3*`data_len]};     
        if (addr == 334) q <= {d[476*`data_len +: 3*`data_len], d[470*`data_len +: 3*`data_len], d[464*`data_len +: 3*`data_len]};     
        if (addr == 335) q <= {d[506*`data_len +: 3*`data_len], d[500*`data_len +: 3*`data_len], d[494*`data_len +: 3*`data_len]};     
        if (addr == 336) q <= {d[536*`data_len +: 3*`data_len], d[530*`data_len +: 3*`data_len], d[524*`data_len +: 3*`data_len]};
        if (addr == 337) q <= {d[566*`data_len +: 3*`data_len], d[560*`data_len +: 3*`data_len], d[554*`data_len +: 3*`data_len]};     
        if (addr == 338) q <= {d[596*`data_len +: 3*`data_len], d[590*`data_len +: 3*`data_len], d[584*`data_len +: 3*`data_len]};     
        if (addr == 339) q <= {d[626*`data_len +: 3*`data_len], d[620*`data_len +: 3*`data_len], d[614*`data_len +: 3*`data_len]};     
        if (addr == 340) q <= {d[656*`data_len +: 3*`data_len], d[650*`data_len +: 3*`data_len], d[644*`data_len +: 3*`data_len]};     
        if (addr == 341) q <= {d[686*`data_len +: 3*`data_len], d[680*`data_len +: 3*`data_len], d[674*`data_len +: 3*`data_len]};     
        if (addr == 342) q <= {d[716*`data_len +: 3*`data_len], d[710*`data_len +: 3*`data_len], d[704*`data_len +: 3*`data_len]};     
        if (addr == 343) q <= {d[746*`data_len +: 3*`data_len], d[740*`data_len +: 3*`data_len], d[734*`data_len +: 3*`data_len]};     
        if (addr == 344) q <= {d[776*`data_len +: 3*`data_len], d[770*`data_len +: 3*`data_len], d[764*`data_len +: 3*`data_len]};     
        if (addr == 345) q <= {d[806*`data_len +: 3*`data_len], d[800*`data_len +: 3*`data_len], d[794*`data_len +: 3*`data_len]};     
        if (addr == 346) q <= {d[836*`data_len +: 3*`data_len], d[830*`data_len +: 3*`data_len], d[824*`data_len +: 3*`data_len]};     
        if (addr == 347) q <= {d[866*`data_len +: 3*`data_len], d[860*`data_len +: 3*`data_len], d[854*`data_len +: 3*`data_len]};     
        if (addr == 348) q <= {d[896*`data_len +: 3*`data_len], d[890*`data_len +: 3*`data_len], d[884*`data_len +: 3*`data_len]};     
        if (addr == 349) q <= {d[926*`data_len +: 3*`data_len], d[920*`data_len +: 3*`data_len], d[914*`data_len +: 3*`data_len]};     
        if (addr == 350) q <= {d[956*`data_len +: 3*`data_len], d[950*`data_len +: 3*`data_len], d[944*`data_len +: 3*`data_len]};     
        if (addr == 351) q <= {d[27*`data_len +: 3*`data_len], d[21*`data_len +: 3*`data_len], d[15*`data_len +: 3*`data_len]};        
        if (addr == 352) q <= {d[57*`data_len +: 3*`data_len], d[51*`data_len +: 3*`data_len], d[45*`data_len +: 3*`data_len]};        
        if (addr == 353) q <= {d[87*`data_len +: 3*`data_len], d[81*`data_len +: 3*`data_len], d[75*`data_len +: 3*`data_len]};        
        if (addr == 354) q <= {d[117*`data_len +: 3*`data_len], d[111*`data_len +: 3*`data_len], d[105*`data_len +: 3*`data_len]};     
        if (addr == 355) q <= {d[147*`data_len +: 3*`data_len], d[141*`data_len +: 3*`data_len], d[135*`data_len +: 3*`data_len]};     
        if (addr == 356) q <= {d[177*`data_len +: 3*`data_len], d[171*`data_len +: 3*`data_len], d[165*`data_len +: 3*`data_len]};     
        if (addr == 357) q <= {d[207*`data_len +: 3*`data_len], d[201*`data_len +: 3*`data_len], d[195*`data_len +: 3*`data_len]};     
        if (addr == 358) q <= {d[237*`data_len +: 3*`data_len], d[231*`data_len +: 3*`data_len], d[225*`data_len +: 3*`data_len]};     
        if (addr == 359) q <= {d[267*`data_len +: 3*`data_len], d[261*`data_len +: 3*`data_len], d[255*`data_len +: 3*`data_len]};     
        if (addr == 360) q <= {d[297*`data_len +: 3*`data_len], d[291*`data_len +: 3*`data_len], d[285*`data_len +: 3*`data_len]};     
        if (addr == 361) q <= {d[327*`data_len +: 3*`data_len], d[321*`data_len +: 3*`data_len], d[315*`data_len +: 3*`data_len]};     
        if (addr == 362) q <= {d[357*`data_len +: 3*`data_len], d[351*`data_len +: 3*`data_len], d[345*`data_len +: 3*`data_len]};     
        if (addr == 363) q <= {d[387*`data_len +: 3*`data_len], d[381*`data_len +: 3*`data_len], d[375*`data_len +: 3*`data_len]};     
        if (addr == 364) q <= {d[417*`data_len +: 3*`data_len], d[411*`data_len +: 3*`data_len], d[405*`data_len +: 3*`data_len]};     
        if (addr == 365) q <= {d[447*`data_len +: 3*`data_len], d[441*`data_len +: 3*`data_len], d[435*`data_len +: 3*`data_len]};     
        if (addr == 366) q <= {d[477*`data_len +: 3*`data_len], d[471*`data_len +: 3*`data_len], d[465*`data_len +: 3*`data_len]};     
        if (addr == 367) q <= {d[507*`data_len +: 3*`data_len], d[501*`data_len +: 3*`data_len], d[495*`data_len +: 3*`data_len]};     
        if (addr == 368) q <= {d[537*`data_len +: 3*`data_len], d[531*`data_len +: 3*`data_len], d[525*`data_len +: 3*`data_len]};     
        if (addr == 369) q <= {d[567*`data_len +: 3*`data_len], d[561*`data_len +: 3*`data_len], d[555*`data_len +: 3*`data_len]};     
        if (addr == 370) q <= {d[597*`data_len +: 3*`data_len], d[591*`data_len +: 3*`data_len], d[585*`data_len +: 3*`data_len]};     
        if (addr == 371) q <= {d[627*`data_len +: 3*`data_len], d[621*`data_len +: 3*`data_len], d[615*`data_len +: 3*`data_len]};     
        if (addr == 372) q <= {d[657*`data_len +: 3*`data_len], d[651*`data_len +: 3*`data_len], d[645*`data_len +: 3*`data_len]};     
        if (addr == 373) q <= {d[687*`data_len +: 3*`data_len], d[681*`data_len +: 3*`data_len], d[675*`data_len +: 3*`data_len]};     
        if (addr == 374) q <= {d[717*`data_len +: 3*`data_len], d[711*`data_len +: 3*`data_len], d[705*`data_len +: 3*`data_len]};     
        if (addr == 375) q <= {d[747*`data_len +: 3*`data_len], d[741*`data_len +: 3*`data_len], d[735*`data_len +: 3*`data_len]};     
        if (addr == 376) q <= {d[777*`data_len +: 3*`data_len], d[771*`data_len +: 3*`data_len], d[765*`data_len +: 3*`data_len]};     
        if (addr == 377) q <= {d[807*`data_len +: 3*`data_len], d[801*`data_len +: 3*`data_len], d[795*`data_len +: 3*`data_len]};     
        if (addr == 378) q <= {d[837*`data_len +: 3*`data_len], d[831*`data_len +: 3*`data_len], d[825*`data_len +: 3*`data_len]};     
        if (addr == 379) q <= {d[867*`data_len +: 3*`data_len], d[861*`data_len +: 3*`data_len], d[855*`data_len +: 3*`data_len]};     
        if (addr == 380) q <= {d[897*`data_len +: 3*`data_len], d[891*`data_len +: 3*`data_len], d[885*`data_len +: 3*`data_len]};     
        if (addr == 381) q <= {d[927*`data_len +: 3*`data_len], d[921*`data_len +: 3*`data_len], d[915*`data_len +: 3*`data_len]};     
        if (addr == 382) q <= {d[957*`data_len +: 3*`data_len], d[951*`data_len +: 3*`data_len], d[945*`data_len +: 3*`data_len]};     
        if (addr == 383) valid <= 1;
      end
    end
    else begin
      init <= 1;
      valid <= 0;
      addr <= 0;
      q <= 0;
    end
  end
  
endmodule