`include "num_data.v"

module w_rom_9 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000000010101000000000001111100000000000100111100111111111110100110111111111100111101000000000000011000111111110010111100111111110101110111000000000011001100;
    mem[1] = 162'b111111111100101010111111111011110011111111111010111000111111111010100001000000000110110011000000000000110010000000000010110110111111111001000000111111111110011110;
    mem[2] = 162'b111111111110000100000000000010011100111111111010110000000000000000011001111111111000111110000000001001101000000000000001000011111111111110001100111111111111111100;
    mem[3] = 162'b111111110100101100111111111001000001000000000000001011111111110011110010111111011111100000000000000111000110000000001000101101111111101001010100111111111100011111;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b000000001010100011111111111011110010111111111000000010111111111111100111000000000000101000111111111110110010000000000100010101000000000100100011000000000011101100;
    mem[33] = 162'b000000000000110000111111111011111001000000000001010100000000000000010001111111111101010111000000000100011001000000000100101111000000000001101111111111110111101001;
    mem[34] = 162'b111111111110011001111111111111110101000000000001100110000000000010111100000000000011100101111111111111110001000000000010001110111111111111111000000000000110101011;
    mem[35] = 162'b111111111110111001000000000100001000000000000000010011000000000010100010111111111101010100000000000000000001111111111010101000111111111010110010000000000110001001;
    mem[36] = 162'b111111111110011010000000000011101101000000000110111010000000000001100110000000000100011101000000000001001101111111111100100000111111110110010001111111111000001001;
    mem[37] = 162'b111111111010011101000000000000111000111111111110010011111111111011110110000000001000101110111111111101011101000000000101010110111111110101101010111111111100110010;
    mem[38] = 162'b000000000010100100000000000011000000000000000101000011000000000010001110000000000010100101000000000001001000000000000011011000111111111110010010111111110110001100;
    mem[39] = 162'b111111111110101100111111111101101111111111111111101100000000000101101010111111111110001111111111111010110011111111111011101001000000000100011001000000000111010111;
    mem[40] = 162'b000000000111101111000000000111001101000000000011100101000000000001000101000000000001001101111111111111110001000000000010100000111111111011111000000000000101110101;
    mem[41] = 162'b000000000101110101000000000001011010111111110111010110000000000001100010000000000101100110111111111100010000111111111101000100111111111011001001000000000000010001;
    mem[42] = 162'b000000000101101000000000000001001101000000000010001101000000000100110011111111111110110001111111111111111011000000000001010010000000000100101010000000000101101000;
    mem[43] = 162'b111111111100011111000000000110010001000000000111110011000000000000100111000000000101000001000000000000000001111111111001111011111111100111100110111111110010101000;
    mem[44] = 162'b000000000101001001111111111111001010111111111111101001000000000000110001000000000010011110000000000100010110111111111001000101000000000010001010000000000011100111;
    mem[45] = 162'b111111111101100100000000001000011101111111111010001110111111111011110001000000000001011101111111111110111100000000000000110110111111111011011001111111111000111010;
    mem[46] = 162'b000000000011110011000000000000011001000000000000010011000000000010110101000000000001000101000000000001111111000000000011000111000000000010011010000000000001111000;
    mem[47] = 162'b111111111111101100111111111011000000111111111111110000000000000110111111111111111010111010111111111110001101000000000011100111000000000011011001000000000100000011;
    mem[48] = 162'b000000000001110011000000000000000100111111111110011010000000000000100101111111111110111010000000000101111110000000001000110011111111111100101111111111111111101100;
    mem[49] = 162'b111111111010001100000000000001100110000000000010010011000000000010101001000000000010110001111111111101101000000000000110011010000000000100000000000000000101101011;
    mem[50] = 162'b000000000011001101000000000110001010000000000011101010111111111001111111000000000000011100000000000001100111111111111101101010000000000010010010000000000101110011;
    mem[51] = 162'b000000000110001101000000001011100001000000000011111001000000000101000111111111111111101011111111111111111110111111111111010101000000000011000101111111111101100000;
    mem[52] = 162'b000000000011001010000000000110000100000000000000011101000000000000001101000000000011101111000000000111101101111111111101110110111111111011110110111111110101010101;
    mem[53] = 162'b000000000101001101111111111001101111111111111100110001111111111101000100000000000010001000000000000101100001000000000001111011111111111101101100000000000100110010;
    mem[54] = 162'b111111111010011100000000000011100011111111111010101001111111111110111110000000000010110111000000000000010001000000000101011011000000000110001110000000000101111111;
    mem[55] = 162'b111111111001001010000000001011011111000000000100101010111111111100101100111111111110111001000000000000000111111111111101000011000000000001111110000000000100101111;
    mem[56] = 162'b111111111000101100000000000100001101111111111111010001111111111111101110000000000000100111111111111011000001000000000000111111111111111110001000000000000000011101;
    mem[57] = 162'b111111111110000100111111111011001010000000000000111011111111111101010000111111111110001111111111111110100110111111111100000111000000000110011011000000000111001000;
    mem[58] = 162'b000000000010001000000000000100100011000000000111100101111111111011100011111111111111001001000000000011111101000000000001111010111111111001010111111111110000010101;
    mem[59] = 162'b111111111011100001111111111111100001000000000000010010111111111111001111111111111101001000000000001000110011000000000000000010000000000001110001111111111000100110;
    mem[60] = 162'b000000000000111110000000000000011000000000000010000101000000000001001010000000000011111100000000000001110101111111111011110111000000000010010111000000000101110101;
    mem[61] = 162'b111111111111100100111111111010101101000000000010010010111111111111110100000000000001000111000000000010001101000000000100101001111111111110001111000000000100101000;
    mem[62] = 162'b000000000010001111111111111111101100000000000101111000111111111100110110000000000000111111000000000011110010111111111101110110000000000000110001000000000100110001;
    mem[63] = 162'b000000000010110101000000000111010000000000000001111101111111111100010101000000000011101001000000000010011100000000000100000010000000000010000110111111111011000101;
    mem[64] = 162'b111111111010111110111111111010110010000000000100101001111111111110011001000000000001001111111111111000101001000000000000000111111111111111101001000000000010010001;
    mem[65] = 162'b111111111110010000000000000010110001000000000010101010111111111110010101000000000001000111111111111010011000111111111010110001000000000101100101000000001001000111;
    mem[66] = 162'b000000001000000001111111111101110110000000000001011001111111110110001100111111111110011100111111111001100100111111111110101110000000000000010101000000000000110011;
    mem[67] = 162'b111111111100110000000000000000000111111111111100000110111111111001111000111111111111010011000000000110111101000000000001010010111111111110001111000000000000000100;
    mem[68] = 162'b111111111101111101000000000000010010000000000001000100111111110111101101000000000010100000000000000001110011000000000001110000111111111011100000111111111110101100;
    mem[69] = 162'b000000000000011100111111111110111100111111111111111101000000000011010101111111111101100011000000000000011101000000000101000100111111111110100100111111111101110101;
    mem[70] = 162'b000000000000000100000000000101110011111111111110011100000000000001111010111111111110001011000000000010110101000000000010011011000000000001001001000000000000000110;
    mem[71] = 162'b111111111011110011000000000001000000111111111100011001111111111111100001111111111111001001000000000000101100000000000011000100000000000101101001111111111101100101;
    mem[72] = 162'b000000000010110000000000000000010011000000000000010101000000000011010010000000000001100101111111111110001011111111111101001110000000000001101100111111111100011001;
    mem[73] = 162'b000000000000000111000000000101001010000000000000101110000000000000111010111111111111001100111111111111010110000000000101010001111111111011010111111111111011001100;
    mem[74] = 162'b000000000100011010111111111111101001000000000001010100000000000010111110111111111110111100111111111111111010000000000110111011000000000011110011000000000010001010;
    mem[75] = 162'b111111111100011001000000000011111001000000000101110111111111111111001011000000000000010000111111111111110011111111111100101111111111111110100001000000000000010110;
    mem[76] = 162'b000000000001011010000000000011000111000000000010101100111111111111110111000000000011001101000000000000010100000000000100000010000000000101110100000000000101000100;
    mem[77] = 162'b111111111110100111111111111101111110111111111100000011000000000010100010000000000000001111000000000101011010000000000100100110111111111101101100000000000100001000;
    mem[78] = 162'b111111111110001000000000000010111000000000000100111001000000000010101101000000000111010111000000000011101001000000000101010101000000000111001100000000000100101011;
    mem[79] = 162'b111111111111011101111111111011011010000000000010101100000000000100111111111111111111100100111111111110010100000000001000000000000000001010000000111111111101101101;
    mem[80] = 162'b000000000011000111000000000010001110000000000001001101111111111101010101111111111101001000111111111111101101000000000001100011111111111101011100111111111011111000;
    mem[81] = 162'b000000000001011011000000000001110100111111111011110101000000000100010111111111111111010111000000000000011010000000000000111010111111111100011010000000001001001000;
    mem[82] = 162'b000000000011001111111111111111010010000000000100001000111111111100110000111111111110000000111111111001000111000000000100111101000000000011001010000000001000100111;
    mem[83] = 162'b111111111111000110000000000100100011000000000101000101111111111100111111000000000000010011000000000001001010000000000001110011000000000110001110000000000000001011;
    mem[84] = 162'b000000000010101011111111111110110000111111111100000111000000000000101001000000000011110110111111110110101010111111111111000100111111111011001100111111111001111001;
    mem[85] = 162'b111111111011010110111111111100000000111111111110001010000000000100001001111111111011010101111111111111111001000000000000000100000000000011010101111111111111111000;
    mem[86] = 162'b000000001000001010000000000100011111000000000000011111000000000100001010000000000001100101000000000001110100000000001000011011000000001000001000000000000110000100;
    mem[87] = 162'b000000000010100101111111111100001011000000000011000000111111111010101110111111111100011101000000000000010000000000000100011001111111111101111100111111111111010110;
    mem[88] = 162'b000000000001100010000000000001100011000000000010011011000000000010001110111111111101101000111111111101010011111111111101010110111111111111101000000000000001010100;
    mem[89] = 162'b000000000000100011000000000000001010111111111101100110000000000001111100111111111110100001000000000000011111000000000010011001111111111110010011111111111000100111;
    mem[90] = 162'b111111111111000110111111111101110011000000000001000110000000000010000010000000000101010010000000000011000001111111111100110011000000000001100110111111111100010000;
    mem[91] = 162'b111111111011010011000000000101010101111111111000100001111111111110100100111111111111000101000000000010101110000000000111001110000000000101000110000000000101011100;
    mem[92] = 162'b111111110110110000111111111111011011111111111100100111000000000000000111111111111111010101000000000010001110111111111001101000111111111101110001111111111000100100;
    mem[93] = 162'b111111111011001110000000000100010001111111111011110000000000000010001000111111111101100110111111111101101101111111111101111000111111111010111010000000000010111101;
    mem[94] = 162'b111111111101001101111111111110100001000000000011000111000000000001001111000000000010011001000000000001001101000000000011010100111111110111010101111111111110110001;
    mem[95] = 162'b111111111111000000000000000011100101111111111111011100000000000100000011111111111101110010000000000100110100000000000110101110111111111110011011111111111100100111;
    mem[96] = 162'b111111111111111001111111111111110000000000000000000100000000000000001100111111111111111000000000000000001011111111111111101111111111111111110100111111111111110101;
    mem[97] = 162'b000000000000001011111111111111110111000000000000010001000000000000000100000000000000001000000000000000000110000000000000001100111111111111111001111111111111111010;
    mem[98] = 162'b111111111111100001111111111111110011111111111111111100111111111111110110000000000000000000111111111111110111000000000000011001000000000000000101000000000000001001;
    mem[99] = 162'b111111111111110100111111111111100110111111111111101110000000000000001001000000000000001000111111111111110000111111111111111001000000000000001110111111111111110011;
    mem[100] = 162'b000000000000001101111111111111111100000000000000000110000000000000001001000000000000000101000000000000001001000000000000000010000000000000000110111111111111111101;
    mem[101] = 162'b000000000000010001111111111111111011111111111111111111111111111111111101000000000000001001111111111111111000111111111111110100111111111111110011111111111111110000;
    mem[102] = 162'b000000000000001010000000000000010011000000000000000101111111111111101010000000000000000011111111111111111101111111111111111111111111111111111111000000000000001000;
    mem[103] = 162'b111111111111111000000000000000011100000000000000001110111111111111111110000000000000001000111111111111111101000000000000000110111111111111110000111111111111101111;
    mem[104] = 162'b111111111111111000111111111111110011000000000000000000111111111111111111111111111111111001111111111111111001000000000000001010000000000000000100000000000000000000;
    mem[105] = 162'b111111111111110110111111111111111011111111111111111101000000000000001001111111111111111000000000000000001000111111111111111011111111111111110011111111111111110101;
    mem[106] = 162'b111111111111111001111111111111111111111111111111111110111111111111111010111111111111110100000000000000000101111111111111111011111111111111101110111111111111110011;
    mem[107] = 162'b000000000000000111111111111111111000111111111111111010111111111111110011111111111111110011111111111111110000111111111111101111111111111111101110000000000000000010;
    mem[108] = 162'b000000000000000110111111111111111100000000000000010111000000000000001110111111111111111111111111111111101111000000000000010110111111111111101011111111111111111010;
    mem[109] = 162'b000000000000000011111111111111101100111111111111110010111111111111111000111111111111111100111111111111111100111111111111101111000000000000000001111111111111111110;
    mem[110] = 162'b111111111111110100000000000000000101111111111111110000111111111111111101000000000000000000111111111111110010000000000000000011111111111111110111000000000000000110;
    mem[111] = 162'b111111111111110111111111111111101101111111111111101010111111111111111001111111111111111101111111111111111001111111111111101010111111111111101101111111111111111010;
    mem[112] = 162'b000000000000010110000000000000010000000000000000110001000000000000001100111111111111010010000000000000010010000000000000011111000000000000000000000000000000110111;
    mem[113] = 162'b000000000000011001000000000000010001000000000000001011000000000000001010000000000000010001000000000000010110000000000000010101000000000000001000000000000000000111;
    mem[114] = 162'b111111111111101010000000000000000010000000000000000000000000000000000101000000000000001001000000000000000100111111111111111011111111111111110100111111111111110011;
    mem[115] = 162'b000000000000001101111111111111101010111111111111111010111111111111111000000000000000000111111111111111110110000000000000001110000000000000000011111111111111111110;
    mem[116] = 162'b000000000000010001000000000000001011111111111111110011000000000000001100000000000000000011111111111111111110000000000000001100000000000000001100000000000000001110;
    mem[117] = 162'b111111111111101111111111111111111010111111111111101011111111111111111101111111111111101111111111111111111001111111111111110100111111111111110110000000000000000101;
    mem[118] = 162'b000000000000000111111111111111111110000000000000000011111111111111111110000000000000000011000000000000011101111111111111111100111111111111110000000000000000000000;
    mem[119] = 162'b000000000000011011000000000000000011000000000000010010000000000000000110000000000000010001000000000000010000000000000000001110000000000000001111000000000000010000;
    mem[120] = 162'b111111111111110100000000000000000001111111111111111001000000000000001101111111111111110101111111111111110010000000000000001001000000000000010011000000000000001101;
    mem[121] = 162'b000000000000000111111111111111111110111111111111011010000000000000001011111111111111111100111111111111111001111111111111111111000000000000000010111111111111111000;
    mem[122] = 162'b111111111111110101000000000000010000111111111111111111111111111111111010111111111111111100111111111111111110111111111111111110000000000000001011000000000000000111;
    mem[123] = 162'b000000000000000000000000000000001000111111111111111011111111111111110110111111111111111110000000000000000101000000000000000000000000000000001001000000000000000000;
    mem[124] = 162'b000000000000000110111111111111111101000000000000001010000000000000001000000000000000000100000000000000000110111111111111111011111111111111111011111111111111111100;
    mem[125] = 162'b111111111111111100000000000000000001111111111111110111111111111111110010111111111111101111111111111111111000111111111111111111111111111111110110000000000000000000;
    mem[126] = 162'b111111111111111101000000000000001111111111111111110100111111111111101101111111111111111010111111111111110101111111111111100111111111111111110001000000000000001011;
    mem[127] = 162'b111111111111111100111111111111111001000000000000010100111111111111111000111111111111110100000000000000011110000000000000000100111111111111111011000000000000000001;
    mem[128] = 162'b000000000000010010000000000010111010111111111110100010111111111111100011111111111111001011000000000000000011000000000001110010111111111111110010111111111111000001;
    mem[129] = 162'b000000000000000011000000000000000010000000000000000010111111111111111110000000000000000000000000000000000110000000000001011001111111111110011111000000000000000010;
    mem[130] = 162'b111111111111110100000000000000000000111111111111111010000000000000000011000000000000000010111111111111111111111111111111111100000000000000000100000000000000000100;
    mem[131] = 162'b000000000000001001111111111111111100000000000000000000000000000000000010000000000000001010000000000000000101111111111111111101111111111111111110111111111111111110;
    mem[132] = 162'b000000000011011010000000000000101111000000000011111111000000000100110110000000000101111011000000000001100000000000000000010101111111111111100100111111111110101000;
    mem[133] = 162'b000000000000000001111111111111110111000000000000000010000000000000000000111111111111111010111111111111111011000000000000000001000000000100100101000000000101000110;
    mem[134] = 162'b000000000000001100111111111111011011111111111111100000111111111111111011000000000000000110000000000000000001000000000000000000000000000000000111111111111111111110;
    mem[135] = 162'b000000000000101010111111111111011101111111111111111001111111111111100101000000000100010010111111111111111000111111111111111011000000000000011001111111111111110111;
    mem[136] = 162'b000000000001010101111111111110001111000000000001010000111111111111010010111111111111110001111111111110101100000000000000001011111111111110110001000000000010000010;
    mem[137] = 162'b111111111111111011111111111111110110000000000000000010111111111111110110111111111111111010111111111111110011000000000010011110000000000011010000000000000101001110;
    mem[138] = 162'b111111111111101111000000000000010111111111111111100001000000000000000001000000000000000111000000000000001000111111111111111010000000000000000000111111111111111011;
    mem[139] = 162'b000000000000100101111111111110111100000000000000000000000000000000000100000000000000000100000000000000000101000000000000101110111111111111111101000000000001110100;
    mem[140] = 162'b111111111111111000111111111111111000000000000000000100000000000000000100000000000000000001000000000000000010111111111111111011000000000000000010000000000000000111;
    mem[141] = 162'b000000000000000011000000000000000000111111111111111011111111111111111001000000000000000011000000000000000011000000000000000101111111111111110011111111111111111101;
    mem[142] = 162'b111111111111111100000000000000000001000000000000000011111111111111111011111111111111111111111111111111111110111111111111111011000000000000000001111111111111111011;
    mem[143] = 162'b111111111111111010000000000000000010111111111111111011000000000000001000000000000000000111111111111111111111000000000000000011000000000000000010111111111111111001;
    mem[144] = 162'b111111111111111111000000000000000100111111111111111111000000000000000001111111111111111100000000000000000001000000000000000001000000000000000010111111111111110111;
    mem[145] = 162'b000000000000000000111111111111111100000000000000000010111111111111111100000000000000000010000000000000000101111111111111111101111111111111111101111111111111111010;
    mem[146] = 162'b111111111111111010000000000000000101111111111111111110000000000000010001111111111111110111000000000000000111000000000000001110111111111111111101000000000000000111;
    mem[147] = 162'b000000000000001110111111111111110010000000000000000101111111111111111000111111111111111010000000000000000101111111111111111111000000000000000010000000000000000001;
    mem[148] = 162'b111111111111110111000000000000000101000000000000000011111111111111111101000000000000000011000000000000000000000000000000000101000000000000000010111111111111111111;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111111111111111110000000000000000011;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule