`include "num_data.v"

module w_rom_21 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b111111111110111001111111111110010000000000000010001011111111111110010001111111111100110001111111111111011111111111110101011000000000000011010100000000000111110101;
    mem[1] = 162'b000000001011000010000000000000011000111111101111000100111111111000100100000000000011111010000000000100110010111111111010101001111111111000011111111111111101100111;
    mem[2] = 162'b000000000010111111111111111100100011000000000001110111000000000001101100111111111110010111111111111110001101111111111111001100000000000001010101000000000100010101;
    mem[3] = 162'b111111101001000100111111101111011000000000000000100101000000010101001100000000010111100110111111110110110100000000000001100011111111101100100101111111111011011001;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111011010010000000000000000100111111111100010101000000000001111111111111111010101011111111110101001011000000000011000111000000000001100100000000000001010000;
    mem[33] = 162'b111111111010000011000000000100000111111111111101010000111111111011000000111111111100010010111111111011001001111111111101100111111111110111101000000000000011010011;
    mem[34] = 162'b000000000010000111000000000010100000111111111001111000111111111101110100111111111011010010000000000000001101000000001000001000000000000000111011111111111111010011;
    mem[35] = 162'b111111111010010001000000000001101111000000000101011010000000000001000000111111111101010111000000000100000100000000000011100100111111111111101010000000001010010001;
    mem[36] = 162'b111111111010010000000000000011001110000000000010101110111111111101110110000000000100110000000000000100111010000000001010001011111111111101010110000000000000110111;
    mem[37] = 162'b000000000011000000111111111101100111111111111011011000111111111001110111111111111111111001111111111111100100111111111100001111111111111111000110000000000101110110;
    mem[38] = 162'b000000000000000110000000000001111011000000000010101000000000000101101001000000000010111110000000001000110011000000000101111111000000000111001011000000000111010101;
    mem[39] = 162'b111111111000101101000000000010110111111111111100110011111111111000100001111111111101000110000000000100000100111111110111110110111111111111100011000000001000011110;
    mem[40] = 162'b000000001000110010000000000010011100000000001000101111000000000000011000111111111011100010000000000100101010000000000000111001000000000100011101000000000010110001;
    mem[41] = 162'b111111111101110010111111111010101100000000000011110011111111110011100001000000001000110001000000000100000001111111111100000100000000000010100100000000000100010111;
    mem[42] = 162'b000000001101001001111111111101010101000000000100001011111111111101110011111111111111000111000000000000110000111111111101100111111111111100011101000000000001001000;
    mem[43] = 162'b000000000000100001000000000011111011111111111111000100111111111100010101111111111101100111000000000100011011000000001010010001000000000110110010000000001000010100;
    mem[44] = 162'b000000000010010100111111111110111010000000000001101110000000000011110111111111111011000111000000000001111110111111110111111001111111111010111000111111111100000111;
    mem[45] = 162'b111111110110101011000000000110111111000000000011101110000000000010000101111111110110000011000000000011001101111111111100101111000000000010110010000000000000001001;
    mem[46] = 162'b111111111001011100000000000001010011000000000010110101111111111110111001111111111110001000000000000100011110111111110101111101111111111000011101111111111001000000;
    mem[47] = 162'b111111111011001111111111111100000001111111111100011111111111111101001000000000000000110001000000000111010100111111111100111011000000000001000011111111111001101100;
    mem[48] = 162'b111111111011110011111111111000010010000000000111000110111111111110001000000000000000100110111111111001010101000000000000001101111111111110011000000000001001101000;
    mem[49] = 162'b000000000101000011111111111010111001111111110111001110111111111101000011000000000000101100000000000101111101111111111110000011111111111010101100111111110110011110;
    mem[50] = 162'b111111111100110000000000000001011000111111111111001110111111111110100001111111111001000110000000000011111010000000001100110011111111111011011100111111111100110101;
    mem[51] = 162'b000000000100101011000000001000011011000000001101110010000000000001010111000000000101110101000000001011110010000000000111000011000000000110011110000000000110011000;
    mem[52] = 162'b000000000010000000000000000011101010000000000100010011000000000101011100000000000101011101000000000101110011000000001001101110000000000000110010000000001110001010;
    mem[53] = 162'b111111111111110101000000000010011100111111111111110011000000000001001010111111111111110101000000000011011011111111111001100111111111111011001110000000000110111001;
    mem[54] = 162'b111111111111100011111111111100010100111111111111110000111111111011000010000000001000001011111111111000111100000000000101010111000000000100101011000000000110101111;
    mem[55] = 162'b111111111011110001000000000010000100000000000010101000000000000101010100111111111011100010111111111101010110000000000110011001000000000010000010111111111100110110;
    mem[56] = 162'b111111111100011100111111110111100111000000000000100111000000000000100100000000000101000011111111111100111000000000000100111000111111110100110010000000000111000001;
    mem[57] = 162'b111111111001000000000000000001100101111111111100110100000000000100100000000000000000101011111111111100111010111111111111101000111111111111011011000000000000000011;
    mem[58] = 162'b111111111101001000000000000001000100000000000001110111000000001101101000000000000001100110111111111101100010000000000100010000000000001000101011000000000010010101;
    mem[59] = 162'b111111111111100110111111111100001001000000000000011010000000000100001110111111111110111111111111111100111001111111111111111010000000000101000100111111111010101111;
    mem[60] = 162'b000000000011111011111111111011010001000000000001001000000000000011010001111111111011100100000000000000110101000000000000010110111111111110101010111111111001001001;
    mem[61] = 162'b111111110110111110000000000010001110111111111110101000000000000000110001000000000010100001000000000100001100000000000000001001111111111100001111111111111011100000;
    mem[62] = 162'b000000000000001100000000000000001010000000000001001001000000000101010011000000000011100101111111111101001111111111111100000111111111111100010101111111111111111111;
    mem[63] = 162'b111111111110110110000000000001110110000000000001000110000000000001010110000000000100010100000000000001001000111111111100100100000000000001101000000000000000100010;
    mem[64] = 162'b111111111011101011000000000001110000000000000000010110111111111110100101000000000100101111000000000011100101000000000000111010000000000011110100111111111111110101;
    mem[65] = 162'b000000000010101110111111111111110000111111111110110001000000000110000011111111111010100100111111111000100111000000000110100100000000000101010011000000000000101010;
    mem[66] = 162'b000000000100001111111111111110001001111111110111100100000000000100111100000000000001010001111111110100010011000000000001111101000000000001101011111111111111110001;
    mem[67] = 162'b111111111100110000111111111010010010111111111110111010000000000001001100000000000010010111000000000001000110111111111100001001000000000000110101000000000011101110;
    mem[68] = 162'b111111111010011110111111111111110101000000000001100111111111111100011010111111111110001100111111111011011110111111111101010100111111111101111000000000000001000110;
    mem[69] = 162'b111111111110101111000000000001001011111111111010011010000000000000101000000000000110111110000000000110000000111111111101011100111111111111100001111111111111001110;
    mem[70] = 162'b000000000000001010000000000000000000111111111100000010111111111000101100000000000010000010000000000010001100000000000000001000111111111111001110000000000000100001;
    mem[71] = 162'b000000000010100011000000000000110010000000000000101111000000000011011011111111111111010111111111111001101001000000000001010110000000000001010000000000000010110010;
    mem[72] = 162'b111111111100110100111111111111110100111111111110110110111111111000000000111111111101111000111111111000100010111111111100101000000000000001100010111111111001001010;
    mem[73] = 162'b111111111011111111111111110110111111000000000001101001000000000001011000000000000100001100000000000000011110000000000001100010000000000001100101111111111100110000;
    mem[74] = 162'b111111111111110110000000000011000110111111110110110111111111111011110010000000000010110101111111111000000101111111111010011011111111111011111110111111111100001001;
    mem[75] = 162'b111111111110010110111111111110110001000000000000101001111111111010110100111111111011010000111111111010100001000000000010110101000000000010110010000000000011010011;
    mem[76] = 162'b000000000100100110000000000111111010000000000001100000000000001010100100000000000100101001000000000000001111000000000111000011000000000011001000000000000111001100;
    mem[77] = 162'b000000000100000010111111111111110011111111111100001101111111111011100011111111111101110100111111111000110011111111110110100101000000000110010011000000000001111000;
    mem[78] = 162'b000000000001001010000000000100100101000000000000100111000000000111111001000000000100001000000000000011110010000000001000110010000000000101010110000000000111110111;
    mem[79] = 162'b000000000011101010000000000011110100000000000010000000111111111010000101000000000100101001111111111101010010000000000010010110111111111111100010000000000011101111;
    mem[80] = 162'b111111111110111000000000000100110011000000000000001001000000000001000011000000000011010001111111111100111001000000000000100001000000000000100010000000000000101111;
    mem[81] = 162'b000000000000010100111111111110000101000000000001011000111111111011111001111111111011000001000000000011111111111111111001110000000000000100110011000000000010110000;
    mem[82] = 162'b000000000000111010111111111111000100111111111111011010000000000001111100000000000010101101000000000000110111000000000010101110111111111001000110111111111110011011;
    mem[83] = 162'b000000000001010100111111111100001011000000000110100001000000000000110010111111111111100111000000000010110011111111111101100101000000000001011001111111111111000111;
    mem[84] = 162'b000000000010000011000000000010000000111111111111010101000000000001101000000000000001110111000000000011110111000000000100000011000000000011100001111111111101110001;
    mem[85] = 162'b000000000001001111111111111111000110111111111100101000000000000110010100000000000000110000000000000111010000000000000000110011000000000101011100000000000000000111;
    mem[86] = 162'b000000000110110000000000000000111100000000000110111011000000000000111111000000000100111101000000001010010100000000000101100000000000001000011001000000000110001101;
    mem[87] = 162'b111111111100011100111111111010101010111111111001001100000000000001111101111111111001101001000000000001001010111111111100000001111111111100100011000000000011000101;
    mem[88] = 162'b111111111001101011000000000000001000000000000011111100111111111110011000000000000001100010000000000010101101111111111010010111111111111010101000111111111111101001;
    mem[89] = 162'b111111111110101110000000000011100110111111111110111110111111111110010100111111111001110010111111111100000100111111111111001011111111111010000000111111111011101010;
    mem[90] = 162'b111111111010100001000000000011001001000000000001110110000000000000110000000000000000111100000000000001000111000000000001011000000000000011110000000000000110110001;
    mem[91] = 162'b111111111110010000000000000011101001111111111100010011111111111011000111000000000011111101000000001000000000111111111111011111111111111011011110000000000100010001;
    mem[92] = 162'b000000000111101011111111111111110100111111111010111110111111111100111110000000000001010010111111111010000100111111111001001011000000000001011011000000000110111000;
    mem[93] = 162'b111111111010110100000000000011110011000000000001110110000000000000010001000000000010000010111111111110000100111111111100110110111111111111001010000000000001101100;
    mem[94] = 162'b111111111001110100000000000101110100111111111101000010111111111101000001111111111101000111111111111110010000111111111110000101000000000010011111000000000001011101;
    mem[95] = 162'b000000000001101100111111111001101011111111111011000001000000000101110001111111111110101001111111111110101000000000000101010100000000000100011001000000000011110001;
    mem[96] = 162'b111111111111011010000000000001010011000000000011011011111111111111010100111111111100110011111111111110000000000000000001011001000000000010010001111111111101001100;
    mem[97] = 162'b000000000001111100111111111111000100000000000010110100000000000010100010111111111111011011111111111110001100111111111101010100111111111011110010111111111110100010;
    mem[98] = 162'b000000000010001111111111111110001000000000000011110111111111111110000001111111111111001111000000000010110101000000000000100010111111111111110011000000000000111100;
    mem[99] = 162'b000000000110101110111111111111000100000000000101111110111111111110001000111111111101000101000000000000111011111111111010001001000000000001001111000000000001000111;
    mem[100] = 162'b000000001000001001000000001001110001000000001011001101000000000111100010000000000101000100000000000100011111111111111011000110111111111110100100000000000010100100;
    mem[101] = 162'b000000000100001110000000000010000100111111111111010111111111111100100111111111111111011011000000000001110011111111111111010100111111111110001100000000000000010001;
    mem[102] = 162'b000000000011110110000000000001101110111111111110100001000000000010010110000000000011001111000000000010100111000000000010010000111111111110000110111111111010101010;
    mem[103] = 162'b000000000001101001000000000000111110000000000001000101111111111111100110111111111101001110000000000001000101111111111100111011111111111111101101111111111011101011;
    mem[104] = 162'b000000000000111111000000000000001100000000000100101010000000000001100100111111111111100101000000000000110010000000000000001111000000000000100001111111111011110010;
    mem[105] = 162'b000000000001001010000000000000111101000000000011000010111111111111011010111111111111000001000000000000000101000000000000100000111111111110011000000000000000000100;
    mem[106] = 162'b111111111010111010111111111010011100111111111010110001111111111110111000111111111101101000111111111110011110111111111101010111000000000000011101111111110111101111;
    mem[107] = 162'b111111111111000110111111111101110100111111110111010111111111110010110001000000000010111111111111111100110011111111111100011010111111111111000100111111111100100110;
    mem[108] = 162'b000000000101001111000000000100001101000000000010000111111111111101100100000000000001001111000000000000101101111111111110010101111111111101110001111111111111010000;
    mem[109] = 162'b000000000011001001111111111111001010111111111110101011111111111011111101111111111110001101111111111111100000111111111100111101000000000000011001000000000010010100;
    mem[110] = 162'b000000000000111100111111111111010110000000000011111000111111111001000110000000000001110111111111111110011000111111111110111101000000000000100000000000000001100000;
    mem[111] = 162'b111111111110010000000000000000011111111111111011111110000000000000110100111111111110010111111111111111111101111111111101100011111111111101010000000000000000111110;
    mem[112] = 162'b000000010100011011000000010001110100000000010001001010000000001110000110000000001110010101000000001010111100000000000011101000000000000101011000000000000000101000;
    mem[113] = 162'b000000000001101001000000000100101101111111111110100100111111111110111101111111111101111011000000000001110000111111111110001011000000000000110111111111111101110100;
    mem[114] = 162'b000000000010100111000000000111001010000000001011001111111111111100111101111111111110111101111111111010111101000000000010100101000000000000001101000000000001101110;
    mem[115] = 162'b111111111101111000000000000010101000111111111101001000111111111111101000111111111101011001111111111010010110000000000001101111111111111111100010111111111110010101;
    mem[116] = 162'b000000000001110111000000000000011010000000000100100101111111111110011101000000000001001110111111111111001110000000000010000000111111111111100100111111111100100011;
    mem[117] = 162'b111111111110101000000000000001001011000000000100010000000000000000110000000000000001011110111111111000111100111111111100001000000000000000100011000000000011000100;
    mem[118] = 162'b000000000100101101000000000000110110000000000011000111000000000000101100000000000000010101000000000001100111000000000001111110111111111101111011111111111111011000;
    mem[119] = 162'b111111111101100100000000000000110000000000000001101101111111111111101101111111111100110101111111111110001000111111111100010011111111111110110111000000000001111110;
    mem[120] = 162'b000000000011000000000000000100111011111111111111111111111111111110001010000000000001110110111111111101000001111111111100010010000000000001001010111111111111010111;
    mem[121] = 162'b000000010000010100000000010001010000000000001110010000000000001111100000000000000110111100000000001010100011000000000011011010000000000000100100000000000101110000;
    mem[122] = 162'b111111111111000111000000000001000010000000000000101001111111111100100101111111111110110011111111111110111010000000000000010011111111111011010011111111111111101011;
    mem[123] = 162'b000000000011111100111111111101101100000000000010001100111111111111001111000000000001000100111111111101110011000000000001110011000000000001000000111111111110110100;
    mem[124] = 162'b111111111111010000000000000101100001000000000011110001000000000100010001000000000001101101111111111101010001000000000001010101111111111110011111111111111111001010;
    mem[125] = 162'b000000000001111100111111111110110110000000000000000001000000000010000001000000000001110110111111110110101100000000000011011000111111111101000001111111111011111110;
    mem[126] = 162'b000000000010100010000000000010101000111111111110010100111111111110001000000000000001010100000000000001101111000000000101011101000000000001110000111111111110100111;
    mem[127] = 162'b111111111110011101000000000001110000000000000010100011000000000000110101111111111101001010000000000001011011111111111101101100111111111111011110111111111111101000;
    mem[128] = 162'b000000000000101111000000000100110101000000000101000110000000000011001011000000000000000111111111111111011101111111111111111000111111111111101011000000000000010110;
    mem[129] = 162'b111111111111111101000000000000000001111111111111111100111111111111111001000000000000000001111111111111111101000000000000000011111111111111011100000000000000001111;
    mem[130] = 162'b000000000000000111111111111111111100000000000000000000000000000000000001111111111111111010000000000000001011000000000000000011000000000000000000000000000000000000;
    mem[131] = 162'b000000000000001001000000000000000000111111111111111100000000000000000110111111111111111011000000000000000000000000000000000101111111111111111011000000000000001011;
    mem[132] = 162'b111111111111111111000000000000000011111111111111110000111111111111110101111111111111010001000000000000000000000000000000010110000000000000100111111111111111100101;
    mem[133] = 162'b000000000000000000111111111111111101000000000000000100000000000000000010000000000000000101000000000000000001111111111111101000000000000000101000111111111111100111;
    mem[134] = 162'b000000000101110010000000000100100000000000000101001110111111111111111001111111111111111111000000000000000010000000000000000010000000000000001011111111111111111011;
    mem[135] = 162'b111111111110011101000000000010111011111111111111101110111111111110111101000000000000111011000000000010000010000000000000011000000000000000010111000000000010111011;
    mem[136] = 162'b000000000000001001111111111111111101000000000000000010111111111111111110000000000000000110000000000000000101000000000000000000000000000000001001000000000000000101;
    mem[137] = 162'b000000000000000011000000000000000011000000000000010011000000000000000101000000000000000000000000000000000010000000000000000000000000000000000000000000000000001010;
    mem[138] = 162'b111111111111111111000000000000000011000000000000000100000000000000001101000000000000010100111111111111111110000000000000001011000000000000000000000000000000000010;
    mem[139] = 162'b111111111111111011000000000000000000000000000000001010000000000000000000000000000000001000111111111111111011000000000000000001111111111111111111000000000000000100;
    mem[140] = 162'b000000000011111001000000000010010101000000000011011101000000000001001000000000000000001101000000000000111110000000000000000010000000000000011001111111111101010101;
    mem[141] = 162'b111111111111110111111111111111110011000000000000000000111111111111111010111111111111110111111111111111110010000000000011010110000000000011011000000000000000011010;
    mem[142] = 162'b000000000011110110000000000100010001000000000101100110111111111111111000111111111111101111111111111111110010111111111111110110111111111111110111111111111111111001;
    mem[143] = 162'b000000000001001100000000000000000100000000000000010000111111111111010011111111111111001010000000000001101010111111111111010010000000000000010111000000000000101001;
    mem[144] = 162'b111111111111110010000000000000000110111111111111110110111111111111110100111111111111110100111111111111111101111111111111111101111111111111111111111111111111111111;
    mem[145] = 162'b000000000000000010000000000000000011000000000000000101111111111111111101000000000000000110000000000000000011111111111111101111000000000000000100111111111111111110;
    mem[146] = 162'b000000000000000011000000000000000000000000000000000010000000000000001100000000000000000100000000000000000111000000000000001100000000000000000010000000000000000010;
    mem[147] = 162'b000000000000000111111111111111111101000000000000000000000000000000000111111111111111111111000000000000000010000000000000000101111111111111111110000000000000000111;
    mem[148] = 162'b111111111111111010000000000000000010111111111111111111000000000000000011111111111111111111000000000000000110000000000000000001111111111111111111000000000000000111;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000010000000000000000001;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule