`include "num_data.v"

module w_rom_31 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b111111111001101111000000000110110000000000000001101011000000000010000100111111111100011110000000000001100110000000000110001100111111111111100101000000000000000010;
    mem[1] = 162'b000000000011011101000000000001100101111111111010101100000000000010100000111111110011111110111111110110010010111111111101110100000000000011100001000000000110000001;
    mem[2] = 162'b000000000011110011111111111001100111111111111110011101111111111111011110111111111111111110111111111111011111111111111001000010000000000010001010111111111000011100;
    mem[3] = 162'b111111011001001000111111100110010000111111101100111010111111100101000011111111101010011011111111111010110110111111100100111011111111101010111111111111111011101000;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b000000001001000110111111111010010100000000000110000000111111111000101011111111111100111100000000000000011101111111111101001000111111111110100100000000000100010111;
    mem[33] = 162'b000000000101110001111111111011011100111111111011111010111111111101111111111111111110100001111111111101000111111111111100011101000000000101110010111111110110011110;
    mem[34] = 162'b000000000100101100111111111010111011111111110110111001000000000100100101000000000101010001111111111101100001111111110110010101111111110001101011000000000101101111;
    mem[35] = 162'b000000000100110100111111111110010011111111111011111100111111111011000000111111110010010011111111111110111010111111111101000101000000000010000101111111110101111000;
    mem[36] = 162'b000000000011011111000000000011001101000000000101001100000000000110100101000000000101001110000000000111011010111111111000010001111111111011101111000000000100000010;
    mem[37] = 162'b111111111001010110111111111110000010000000000001111011111111111110100010000000000111110111111111111110011001111111111011001110000000000000011000111111110010100000;
    mem[38] = 162'b000000000110110001000000000100001111000000000111010010000000001011000000111111111110111010111111111111100101000000000100100000000000000011100000111111111010101001;
    mem[39] = 162'b000000000000110100000000000001001101111111111010110111000000000010001101000000000010101000111111111000011101111111110110110001111111111100011000000000000010111000;
    mem[40] = 162'b000000000100111000000000000101000010000000000100101101000000000000101111111111111110101011000000001000001111000000000100111010000000000010100111000000000010011011;
    mem[41] = 162'b111111111100110001111111111110001110000000000110111101111111111010100110000000000000101101000000001011001100111111111001100001111111111110000011111111111100111110;
    mem[42] = 162'b000000000000001101000000001010100110111111111111111111111111111011110111111111111011111001000000000010100101111111111100000100111111111111100100000000000101101000;
    mem[43] = 162'b000000000011111110000000000001111111000000000100111010000000000110001001111111111001110011000000000100001110000000000101000011111111111010010100111111111011100000;
    mem[44] = 162'b000000000010111000000000000100100011000000000010000010111111111111111101111111111110000001111111111101011111000000000010010000111111111011000101000000000010001010;
    mem[45] = 162'b111111111010000000111111110111100110111111111101001011111111111011111011111111111000101100111111111101011011111111111010111000111111111100100010000000000010001001;
    mem[46] = 162'b111111110110100001000000000011011000111111111111011100111111111101111111111111111110101110111111111011110111000000000010000000111111111010001001000000000001001001;
    mem[47] = 162'b000000000011011101111111111100010011111111110011110001000000000101110001111111110111000010000000000010111100000000000000010000000000000000000101000000000100010000;
    mem[48] = 162'b111111111001111110111111111110101100111111111111010011000000000000100000111111111000110101000000000110110011111111110100111101111111110110100011111111111110110101;
    mem[49] = 162'b111111110100101110111111111010010010111111110111111100000000000010100011000000000110001001000000000011101110000000000000010000000000000110110111111111110110101100;
    mem[50] = 162'b000000000011000100000000000000101000000000000100011010000000000000001111111111111011101011111111111111110010000000001000101000111111111111000110000000000010010001;
    mem[51] = 162'b000000000110010101000000000001000011000000000101000101000000001101101010000000000100101110000000000000100101000000000111101011000000000111011100111111111110101111;
    mem[52] = 162'b000000000110001001000000000001000011000000000000111010000000000100111011111111111101011001000000000001110101000000000111110100111111111111111111000000000100001101;
    mem[53] = 162'b000000000001011011111111110110101010111111111110110001000000000000000010111111111110011100111111111100111000111111111110100010000000000110000001111111111110011001;
    mem[54] = 162'b000000000001110100111111111011111101000000000001000110111111111111110001000000000000101011111111111110100001000000000001000110111111111100101101111111111010111111;
    mem[55] = 162'b000000000101101111111111111101101110000000000111001010111111111101111001111111111011001110111111111101110110000000000011111100000000000000011000000000000001111111;
    mem[56] = 162'b111111111100010111000000000100110011000000000010001100111111110111100001000000000000000100111111111111101000111111111011000000111111111100011100000000000000010010;
    mem[57] = 162'b000000000111001000111111111110011110111111111111010111000000000001101001111111111100011110000000000000011100111111111010100011111111111110111110111111111111101100;
    mem[58] = 162'b000000000010010001000000000001110010000000000101011110111111111111100101111111111111000001000000000000001010000000000100001010111111111111001011111111111010011001;
    mem[59] = 162'b000000000001010110000000000100000111000000000001001010000000000000101100111111111101010110111111111110101000000000000001000001111111111011010001111111111001111110;
    mem[60] = 162'b000000000111111000000000000010000001111111110110100111000000000100000111000000000011111110111111110110010100111111111100111100000000000100111110000000000010010011;
    mem[61] = 162'b000000000001110110000000000011101001111111111011011111000000000011110111000000000001110111000000000000111110000000000001010001000000000111010000111111111110001100;
    mem[62] = 162'b111111111010101000000000000001101111000000001000010111111111111101101111111111111111001110111111111011111110000000000100011110111111111101010000000000001000000101;
    mem[63] = 162'b111111111110111110000000000100100000000000000011100010000000000011011101000000000101101111000000000010010000000000000101111001111111111100111110111111111011100101;
    mem[64] = 162'b000000000100100010111111111101111111111111111010011110111111111010110100000000000000101100111111111110101011000000000001010000000000000001010001111111111110110011;
    mem[65] = 162'b111111110110110010111111111110110111111111111111001000111111111101001110000000000000110101000000000000000101000000000010001110000000000110011011000000000001000000;
    mem[66] = 162'b111111111101000010000000000010001110111111111001011011000000000100100111000000000000111100000000000001111111111111111011110111111111111111100101111111111101110011;
    mem[67] = 162'b111111111110101011111111111110000011111111111010111001111111111101101010111111111010010101111111111010011100000000000001110011111111111111101010000000000000000001;
    mem[68] = 162'b111111111110001101111111111101000111111111111001111101111111111110001100000000000010011111000000000010111101000000000010010111000000000000000010111111111001101000;
    mem[69] = 162'b000000000000101100111111111100110110111111111101111011000000000000010010000000000100001101000000000001111010000000000001010101000000000100110010000000000001000000;
    mem[70] = 162'b111111111010000010000000000010100111111111111110101101111111111101100010000000000101001101111111111110100110111111111110001100000000000001001100000000000011011110;
    mem[71] = 162'b111111111101011011111111111111010011000000000010010010000000000001110001000000000010001010111111111110011000000000000010011011111111111100011000111111111100000101;
    mem[72] = 162'b000000000000110110111111111101101100111111111000000001111111111000111110111111111111000010111111111011101100000000000000000110111111111111111111111111111100101111;
    mem[73] = 162'b000000000001000100000000000000011010111111111010100101000000000001010010000000000000010101000000000010011100000000000001110011111111111111101000111111111010000011;
    mem[74] = 162'b000000000000101010111111111110111110111111111100111000111111111101100011000000000011000000111111111111000100000000000001001010000000000000011111000000000100100000;
    mem[75] = 162'b111111111001010110111111111110011001111111111110000000000000000001100001000000000011110110111111111111111111111111111011101011000000000010101001000000000100011101;
    mem[76] = 162'b111111111111110100000000000000110011111111111110111101000000000111010000000000000010101001000000000111111100000000000110001010000000000000101011000000000010111011;
    mem[77] = 162'b000000000000100100111111111111101001000000000110100101111111111101111101000000000000101101111111111111101101000000000011100101000000000010011101000000000000111000;
    mem[78] = 162'b000000000001110100000000000000100001000000000100110110000000001000100101000000000111010111000000000100111110000000000011000101111111111111011001000000000101011000;
    mem[79] = 162'b111111111010001010000000000001110001000000000100001001111111111110011001111111111010000110000000000010000000111111111111010011111111111010101110000000000010011011;
    mem[80] = 162'b111111111101011101000000000000011111111111111001000001000000000001111011000000000011100010000000000010001001111111111111000101111111111010110111000000000010011010;
    mem[81] = 162'b111111111110001110111111111100110000111111111111100110111111111010000110111111111101001000000000000101100110000000000001111011111111111011101000000000000100100111;
    mem[82] = 162'b000000000000100111111111111111011111000000000001110000000000000010001011000000000010100011111111111110010100111111111111100011111111111010111111111111111110010101;
    mem[83] = 162'b111111111000110001000000000010011011000000000001101000000000000001111001111111111111001000111111111001000011111111111110001000000000000000100110000000000101101001;
    mem[84] = 162'b111111111010100110111111111111001000000000000010101001111111111011111101000000000100100101111111111100010011111111111011011010111111111101101011000000000001101100;
    mem[85] = 162'b000000000000001011111111111111000111000000000010111100111111111100111010000000000011110100000000000011001100111111111111100000000000000000010010000000000011011011;
    mem[86] = 162'b111111111101011111000000000001010011000000000100100011000000000001001111000000000011001011000000000101110000000000000011100101000000000100111100000000000111110011;
    mem[87] = 162'b000000000000000000111111111101000101111111111110100010111111111111000111111111111100100011111111111111111011111111111101111001111111111010010000000000000001000011;
    mem[88] = 162'b000000000001001101000000000010010001111111111100110101000000000001011110000000000100010001111111111100111101111111111110100100000000000011000010111111111000110010;
    mem[89] = 162'b000000000000110100111111111101001000111111111111000011111111111100101111000000000010111110000000000000101011111111111100101010000000000001000101111111111111100010;
    mem[90] = 162'b000000000101010000000000000101010001000000000000111011111111111111101101111111111101111101111111111111000101111111111111001010000000000011001001000000000011010010;
    mem[91] = 162'b111111111110101100000000000010011110000000000011010001000000000001000010111111111111001010000000000011000101000000000010001001000000000000111001000000000010000000;
    mem[92] = 162'b000000000000100101000000000010110001111111111101011011000000000001111100111111111111011000111111111110010011111111111111011111000000000000010101111111111111111001;
    mem[93] = 162'b000000000100101111000000000000100100111111111001010110111111111110011000111111111010011110000000000011101100111111111111001011000000000110100001111111111100110011;
    mem[94] = 162'b111111111111000001000000000011111000111111111000101111000000000001101100111111111011011001111111111111100001111111111110101101111111111001010001111111110111001100;
    mem[95] = 162'b111111111100001010111111111101000111000000000101011111000000000100001101000000000010010000111111111110111011000000000001111110000000000001101000000000000010000111;
    mem[96] = 162'b000000000000000111111111111111110110000000000000011001000000000000001011000000000000000010000000000000001101111111111111100001111111111111101100000000000000000010;
    mem[97] = 162'b000000000000001100000000000000001000000000000000011000000000000000110011000000000000010101111111111111101101000000000000010000111111111111101011111111111111110101;
    mem[98] = 162'b111111111111110001000000000000000101000000000000000011000000000000100000000000000000100111111111111111111000000000000000100100111111111111110110111111111111111100;
    mem[99] = 162'b000000000000001110000000000000001110000000000000011001111111111111101110000000000000000001000000000000010010111111111111100100111111111111111110111111111111110110;
    mem[100] = 162'b000000000000010111000000000000010000000000000000001100000000000000000001000000000000001011000000000000001011000000000000001000000000000000001010000000000000001111;
    mem[101] = 162'b000000000000010111000000000000000100000000000000100000000000000000001011000000000000001110000000000000000011111111111111111101111111111111111000111111111111111001;
    mem[102] = 162'b111111111111111110111111111111111110111111111111110001111111111111111111000000000000001001000000000000001001000000000000001110000000000000000010000000000000000100;
    mem[103] = 162'b111111111111111010000000000000001001000000000000000111111111111111111010000000000000001111000000000000001110000000000000011010111111111111111100111111111111101111;
    mem[104] = 162'b000000000000010110000000000000010000000000000000001101000000000000011010000000000000001001000000000000010001000000000000011001000000000000010000000000000000001001;
    mem[105] = 162'b111111111111100111111111111111110001000000000000100000000000000000000111111111111111111000000000000000000110000000000000001010000000000000001100111111111111101110;
    mem[106] = 162'b000000000000010010000000000000010100111111111111110010000000000000011011000000000000001101000000000000011101000000000000001000111111111111111100000000000000001110;
    mem[107] = 162'b111111111111101000111111111111101100111111111111111110111111111111110110111111111111110010111111111111101101000000000000010100000000000000010001000000000000010110;
    mem[108] = 162'b000000000000010001000000000000010010000000000000010111000000000000000100111111111111111100000000000000001110000000000000010000000000000000000001111111111111111101;
    mem[109] = 162'b000000000000101010000000000000010000000000000000010000000000000000001111000000000000000110111111111111111111111111111111110111000000000000010011000000000000001001;
    mem[110] = 162'b111111111111111100000000000000010000000000000000000110111111111111110000000000000000000110111111111111111001000000000000010010111111111111111101000000000000000100;
    mem[111] = 162'b000000000000000011000000000000000011000000000000000111000000000000000000111111111111111101000000000000000010111111111111111011000000000000000011000000000000001010;
    mem[112] = 162'b000000000000100010000000000000101101000000000000011010000000000000000101111111111111111010000000000000100110111111111111111001111111111111111100000000000000011111;
    mem[113] = 162'b000000000000011000111111111111111101000000000000000001000000000000000001000000000000000101000000000000001101000000000000000010000000000000000010000000000000010011;
    mem[114] = 162'b000000000000000111000000000000010011111111111111110111111111111111110011111111111111111101000000000000001111111111111111110111111111111111111010000000000000001110;
    mem[115] = 162'b111111111111110001111111111111010110000000000000010010111111111111111011000000000000010100000000000000001000000000000000001001000000000000010101000000000000010011;
    mem[116] = 162'b111111111111111010111111111111110011111111111111110101111111111111001100111111111111101101000000000000000001111111111111111001111111111111110000000000000000000100;
    mem[117] = 162'b000000000000001100000000000000001111111111111111101111000000000000010000111111111111110001111111111111101110000000000000001010000000000000000100000000000000011001;
    mem[118] = 162'b000000000000010000000000000000010010000000000000001001000000000000011000000000000000000011111111111111111001000000000000010110000000000000000011000000000000010001;
    mem[119] = 162'b111111111111111010111111111111110111111111111111110000000000000000000011000000000000001100000000000000001101111111111111111000000000000000000001000000000000001110;
    mem[120] = 162'b000000000000001101000000000000011100000000000000000100000000000000010001000000000000000111000000000000001110000000000000010010000000000000011111000000000000000000;
    mem[121] = 162'b000000000000011100000000000000001001000000000000011101000000000000011011000000000000011001000000000000010101000000000001001011000000000000100000000000000000010110;
    mem[122] = 162'b111111111111111111000000000000011011111111111111111011000000000000001000000000000000000110000000000000000101111111111111110010000000000000001100000000000000010101;
    mem[123] = 162'b111111111111111110000000000000001101000000000000001110000000000000000110000000000000000100111111111111110101111111111111111000111111111111111011111111111111110001;
    mem[124] = 162'b000000000000010001111111111111111111000000000000011010000000000000000001000000000000001010000000000000001101000000000000000100000000000000000010000000000000000110;
    mem[125] = 162'b111111111111101001111111111111110101111111111111101000111111111111110000111111111111111101111111111111111000000000000000100001000000000000011010000000000000011010;
    mem[126] = 162'b000000000000010100000000000000001001111111111111111001111111111111111001111111111111101110111111111111111110000000000000011000000000000000001110000000000000100001;
    mem[127] = 162'b000000000000000111111111111111110010000000000000001111111111111111101011111111111111110011111111111111111011111111111111011100111111111111110000111111111111111100;
    mem[128] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[129] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[130] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[131] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[132] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[133] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[134] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[135] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[136] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[137] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[138] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[139] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[140] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[141] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[142] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[143] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[144] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[145] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[146] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[147] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[148] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule