`include "num_data.v"

module w_rom_1 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b111111111100011000111111111100011001111111111000100110111111111010001001111111111110101101111111111111011010111111111111100011000000000000011010000000000011011101;
    mem[1] = 162'b111111111101111000000000000111111110000000000111010001000000000111100001111111111010011110000000000101110001000000001010100000111111110101100000000000000010101010;
    mem[2] = 162'b000000000010001011111111111111000100000000000001110001000000000001110010000000000000111000000000000010001100000000000010001000111111111111110101111111111010100111;
    mem[3] = 162'b111111100000010001000000000111011010111111111010011000000000000011010111000000011110010101111111110011011001111111110111100010111111110001000000111111110000111101;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111000010111111111111110011000000000000000010101000000000000011010000000000000000111111111111001000000111111111000100110111111111110000010000000000101010001;
    mem[33] = 162'b000000000110010010000000000100001011111111111010001000111111110110100100000000000011100100111111111111111111111111111001000011000000000011001000111111110111111111;
    mem[34] = 162'b111111111100110111111111111010110100000000000001101000111111110111111001000000000000011101000000000010000110111111111111000101111111110110101111000000000011110010;
    mem[35] = 162'b111111111111000000000000000001001111000000000000111000111111111011010111111111111000010111000000000001011110000000001011111000000000000000001011000000000100101110;
    mem[36] = 162'b000000000010000100000000000000001011000000000001010001000000000010101110111111111101010010111111111101110100000000000011001110111111111110100001111111111101000011;
    mem[37] = 162'b000000000001001100111111111110100110000000000001000000000000000000011110000000000110110100111111110111100000000000000010001011111111111000111100111111111000011001;
    mem[38] = 162'b000000000011001000000000000101000110000000000100101001111111111111011010000000000010111110111111111111010011111111111110001110000000000111111100000000000111011100;
    mem[39] = 162'b000000000011011111000000000011110100111111110011100101111111110111011000000000000011111001111111111111011001000000000001011000111111111100111110111111111110001001;
    mem[40] = 162'b000000000100000111000000000000110100000000000110000110000000000000000001111111111101101111000000001010000011000000000000001001111111111001100110000000001111011011;
    mem[41] = 162'b000000000001011001111111110110101111000000000010000110111111111010010000111111111111010111000000000010010011111111111110011001000000000100000111000000000101101101;
    mem[42] = 162'b111111111011000101111111111101101110000000000000010110000000000110100001111111111011000101111111111011010101111111111101010011000000000000000110000000000101100100;
    mem[43] = 162'b000000000110000000000000000100010011000000000011100001000000000011011011000000000000101110000000000000110001000000001000000001000000000100100101000000000111111100;
    mem[44] = 162'b000000000101001100111111111111001111111111111100001000111111111111011101111111111101000011000000000001110101111111111101001010000000001000001100111111111100011111;
    mem[45] = 162'b000000001100001101000000000001011110000000001000010010111111111001001110000000000000100111111111111000010100000000000001011101000000000011000011111111111011000110;
    mem[46] = 162'b000000000001001011000000000100100110000000000111011110111111111101011100111111111000101001000000000011110011111111110001010001000000000110101101000000000000010110;
    mem[47] = 162'b111111111100000101111111110111011000000000001010000001111111111110100001111111110110101011000000000101111101111111111010110000000000000111100110111111111110011001;
    mem[48] = 162'b000000000101010110111111111000000111000000000110100101111111111110011000000000000010101001000000000001000010111111111110010000000000000011000000000000000011000111;
    mem[49] = 162'b000000000011111111000000000010001100000000000010101111111111111101100100000000000111001111000000000000000101111111111110110010111111111101000011111111111100000111;
    mem[50] = 162'b111111111110010100000000000010010000111111111110011111111111111111100101111111111010010010000000000110001010111111111011010111000000000010101000000000000001101111;
    mem[51] = 162'b000000001100000000000000001000010101000000001101000100000000000101000001000000000011010000000000000111011011000000000110000001000000000100010001000000001001001001;
    mem[52] = 162'b000000000000110001000000000110111101000000000100101000000000000100000100000000000000010010000000000010000110000000000101001111000000000011010110000000000010000111;
    mem[53] = 162'b000000000000101010111111111011101000000000000010101101111111111110011100000000000010010011000000000110101000111111110111111000000000000000011010000000000010111110;
    mem[54] = 162'b000000000100101101111111110110101010000000000000000110000000000100111011000000000101011010111111110110111111000000000011001101000000000000000001111111111011100101;
    mem[55] = 162'b111111111001000111000000000000111110111111111101011010000000000001100001111111111000011101111111111110011110111111111100111010000000001001101001000000000011101111;
    mem[56] = 162'b111111110000101001000000001101000111111111110010010101111111111111100100111111111101011111111111111001010110111111110011110111000000000101111000000000000110110101;
    mem[57] = 162'b000000000001101110000000001001111101111111110000001100111111111111001101111111111110010010111111111100101010000000000000010100111111111110111000000000000001110111;
    mem[58] = 162'b000000000011100000000000000001100000111111111111011000000000000000101011000000000011100100111111111110011111000000000111010101000000001010101011111111111110100010;
    mem[59] = 162'b000000000111100000000000000100000010111111111011010100000000000001000000000000000110010111000000000001001010111111111100110100000000000011111111111111110011000100;
    mem[60] = 162'b000000000000110000111111111100101001000000000001011111111111111101010100111111111010000111000000000011110010000000000110110000111111110110110101000000000000100001;
    mem[61] = 162'b000000000010001000111111111100000111000000000100001001000000000000010100000000000001011000000000000100010001111111111111110100000000000011011011111111111101100101;
    mem[62] = 162'b111111111011101000111111111110010011000000000001011101111111111110110110000000000100100010000000000000001110000000000100111100000000000001000001000000001000001010;
    mem[63] = 162'b000000000011010010111111111100000101111111111111111110111111111110010001000000000001111011000000000101001001111111111000001110000000000001100001111111111100011001;
    mem[64] = 162'b111111111111111100111111111101010011000000000100010111111111111110001100000000000100011111000000000000001010000000000000101011000000000001100000111111111101100100;
    mem[65] = 162'b000000000001110101111111111101101111111111111011100100000000000010111000111111111110111111111111111111010000111111111101011000111111111101111001111111111101001101;
    mem[66] = 162'b000000000011011110000000000011010010000000000000101001111111111110010000111111111101100111000000000000110101000000000010011000111111111101110110111111111101101100;
    mem[67] = 162'b000000000010001111000000000000001101111111111111100111000000000001001100111111111111101011111111111101011010000000000000001111111111111011111101111111111000010111;
    mem[68] = 162'b111111111111110101000000000001101101000000000011110010111111111110101101111111111110011000111111111111110000111111111101110010111111111001111100000000000001001011;
    mem[69] = 162'b000000000100001101111111111111110101111111111111110101111111111110011111111111111010111111000000000001100000111111111110110001111111111101001110111111111111100010;
    mem[70] = 162'b000000000101100110111111111101010001111111111110111101111111111010010100000000000000010100000000000110101110111111111100101011111111111111111001111111111111001001;
    mem[71] = 162'b111111111001111100111111111011010011111111111100111101111111111111100100000000000010011001111111111011110101111111111111000100111111111100111001111111111111010111;
    mem[72] = 162'b000000000110000000111111111101010011111111111011101110000000000011000101111111111101001111000000000010001110111111111101010110111111111101011010111111111001111111;
    mem[73] = 162'b111111111110100010000000000001010001111111111100111110000000000010010100000000000000010110000000000000111010000000000000010000000000000000000001111111110110011100;
    mem[74] = 162'b000000000100110000111111111010010101111111111101010001111111111111010101111111111111001100111111111101000010000000000101001111111111111111010111000000000001010000;
    mem[75] = 162'b111111111101110001000000000000010010000000000000000011111111111011010011000000000000011100000000000010000110111111111010100101000000000000110111111111111100110010;
    mem[76] = 162'b000000000110011111000000000010111000111111111101101010000000000100110010000000000010101100000000000100011100000000000010111110000000000111100111000000000101110110;
    mem[77] = 162'b111111111111100010000000000110000010111111111011011010111111111111000110111111111110100010000000000000110011111111111000010110000000000000001111111111111110111100;
    mem[78] = 162'b000000000000100100000000000101110101000000000011110011000000000011100011000000000101111110000000001010010111000000000010001010000000000010100110000000000100100010;
    mem[79] = 162'b111111111011011110000000000001101110111111111110100001111111111111011001111111111100110011111111111110101101000000000110110100000000000000100001000000000011111110;
    mem[80] = 162'b000000001000111101000000000010100110111111111101100001000000000010100000111111111110110011111111111111001010111111111110110111111111111101011001111111111000111001;
    mem[81] = 162'b111111111100010000000000000010000011111111111111001101000000000001001101111111111111110000111111111111111100111111111110010011000000000001100001000000000000110010;
    mem[82] = 162'b111111111111110011000000000010011100000000001000000110000000000001111101000000000000001010000000000100100100111111111001000101000000000000111010111111111011100010;
    mem[83] = 162'b111111111101100101000000000011100000000000000000000011000000000011101011111111111111001101000000000011001101111111111011111101000000000010001110111111111111001001;
    mem[84] = 162'b111111111101101011111111111011000100000000000001000100111111111101111110000000000010110010000000000000000110111111110011101000000000000010010011000000000000111110;
    mem[85] = 162'b000000000000110111111111111111000011000000000010110111111111111111110101000000000010010000000000000000000000000000000000010011000000000100000011111111111110001110;
    mem[86] = 162'b111111111110100110000000000001100010000000000000010001000000000111011100000000000101101001111111111110010010000000000011010101000000000110101110000000000100111000;
    mem[87] = 162'b111111111111010100111111111110000100000000000011111001111111111100100101111111110110100010000000000000101000000000000001111000000000000000011011000000000001111001;
    mem[88] = 162'b000000000010011111111111111111011001111111110110110110111111111101010101000000000010010010111111111011011101111111111000001100000000000000000010000000000110010100;
    mem[89] = 162'b000000000100110100111111111111101011111111111110010000000000000011011110111111111101101001111111111101110010111111111111110000000000000001011010111111111001000010;
    mem[90] = 162'b000000000010111101111111111101100001000000000010010101111111111101011001000000000001100010111111111111001011000000000001011011000000000101101100000000000100111110;
    mem[91] = 162'b000000001000000001000000000000010100000000000100010101000000000010101101111111111100111110111111111111000101000000000011001101000000000010011100000000000100000011;
    mem[92] = 162'b111111111110110110000000000010101111000000000000110001000000000000001100000000000010010001111111111100010110111111111111010111111111111110001110111111111010001001;
    mem[93] = 162'b111111111111101011111111111101100000000000000101110001111111111011101010000000000001001101111111111110100110111111111111110100111111111100001001111111111111001100;
    mem[94] = 162'b111111111110001011000000000001111111000000000010011110000000000010001010111111111101110110111111111110111100000000000000111100000000000000011110111111111010011000;
    mem[95] = 162'b000000000010011111000000000011001001000000000010111101000000001000000110111111111111000100000000000001100010000000000110100000111111111101100110111111111101001010;
    mem[96] = 162'b000000000000001111000000000000001101000000000000001100111111111111111001111111111111111011111111111111110101111111111111100101000000000000000010000000000000001010;
    mem[97] = 162'b000000000000000000000000000000000010000000000000000000111111111111110000111111111111110101111111111111111010000000000000000001000000000000000111000000000000000010;
    mem[98] = 162'b000000000000000001111111111111101011000000000000100000000000000000000111111111111111111010000000000000000100000000000000011110000000000000001011000000000000000111;
    mem[99] = 162'b111111111111100110111111111111111010111111111111101001000000000000001000000000000000000110111111111111111010111111111111111101111111111111110111000000000000000101;
    mem[100] = 162'b111111111111110101000000000000000010111111111111111111000000000000001101111111111111111111000000000000010110000000000000000010111111111111111011000000000000011111;
    mem[101] = 162'b000000000000001100111111111111111110111111111111011100000000000000001110000000000000000001000000000000010101111111111111110101111111111111110100000000000000000001;
    mem[102] = 162'b111111111111110010111111111111111010000000000000001010000000000000001001000000000000001000000000000000000101000000000000001100111111111111111001111111111111110111;
    mem[103] = 162'b111111111111111001000000000000000000000000000000001010111111111111111100000000000000010010000000000000001000000000000000010010000000000000000101000000000000000010;
    mem[104] = 162'b000000000000001001111111111111110111111111111111101000111111111111111001000000000000000110111111111111111011000000000000001111000000000000000110000000000000010101;
    mem[105] = 162'b111111111111110001111111111111111000111111111111111001111111111111111111111111111111111110000000000000000000111111111111111011111111111111111010000000000000001001;
    mem[106] = 162'b111111111111111001111111111111110110111111111111111010111111111111101111111111111111111011000000000000000000000000000000001010111111111111111101111111111111110111;
    mem[107] = 162'b111111111111111111000000000000000010000000000000000001111111111111110011111111111111111100111111111111110100111111111111110001111111111111111000111111111111111110;
    mem[108] = 162'b111111111111110000111111111111111100000000000000001010000000000000001110000000000000001101000000000000001000000000000000000000000000000000000011000000000000001100;
    mem[109] = 162'b111111111111111001111111111111111001000000000000001000111111111111111100111111111111111101111111111111111101000000000000001010111111111111111111111111111111110010;
    mem[110] = 162'b111111111111101011000000000000000111111111111111111010111111111111111001111111111111111001111111111111111101111111111111110111000000000000001100111111111111111110;
    mem[111] = 162'b000000000000010010111111111111110111111111111111100101111111111111110101111111111111111101000000000000001100111111111111100100111111111111111011111111111111110111;
    mem[112] = 162'b000000000000101111000000000000000011000000000000011001000000000000001000111111111111111100111111111111111101000000000001000010000000000000000011000000000000000111;
    mem[113] = 162'b000000000000000101000000000000000101111111111111011011000000000000000001000000000000000110000000000000001000000000000000010010000000000000001011000000000000010010;
    mem[114] = 162'b111111111111111010000000000000000000000000000000001011111111111111111011000000000000000001000000000000000101111111111111111010000000000000001000000000000000001011;
    mem[115] = 162'b111111111111111010000000000000000001000000000000000000111111111111111100111111111111111001111111111111110110000000000000000001000000000000000001000000000000000011;
    mem[116] = 162'b000000000000011001000000000000000000000000000000011101111111111111111011111111111111110001000000000000001010000000000000001110000000000000001011000000000000000001;
    mem[117] = 162'b000000000000001110111111111111110101000000000000010101111111111111011111111111111111110101000000000000000100000000000000001000000000000000000001000000000000000010;
    mem[118] = 162'b111111111111111111000000000000001101000000000000010110111111111111111010000000000000000000000000000000001000111111111111111101000000000000001100000000000000000010;
    mem[119] = 162'b000000000000000000000000000000000000111111111111101111000000000000000001000000000000000011111111111111101111111111111111110011000000000000000111000000000000000111;
    mem[120] = 162'b111111111111101110000000000000000000000000000000010000111111111111101101000000000000000110111111111111110001111111111111111001111111111111111000000000000000000001;
    mem[121] = 162'b000000000000001000000000000000000110111111111111110110000000000000001111111111111111111001000000000000010001111111111111101001111111111111111110000000000000101001;
    mem[122] = 162'b000000000000011101000000000000000000000000000000000000111111111111110111111111111111101101111111111111101110000000000000100100000000000000000011111111111111111110;
    mem[123] = 162'b111111111111111100000000000000001001111111111111110000111111111111111100000000000000000000000000000000000001000000000000000100000000000000000111111111111111111010;
    mem[124] = 162'b111111111111101001111111111111111001111111111111110111000000000000001000000000000000001101111111111111110011000000000000001100111111111111110001111111111111111101;
    mem[125] = 162'b111111111111110111000000000000000001000000000000001011000000000000000000000000000000000010111111111111110111000000000000001101111111111111111111111111111111111100;
    mem[126] = 162'b111111111111110110000000000000001001111111111111100101111111111111111001000000000000000000111111111111100111111111111111111011111111111111111111000000000000000111;
    mem[127] = 162'b000000000000001101000000000000000100000000000000000101000000000000001001000000000000001001000000000000001111111111111111111100000000000000001001000000000000001000;
    mem[128] = 162'b111111111100111001000000000001100111111111111100101011000000000000001111000000000000010011111111111111100000000000000000111000000000000000011001111111111101101000;
    mem[129] = 162'b000000000000000111000000000000000011000000000000000001000000000000000100111111111111111110000000000000000011111111111111110100111111111101110110000000000001000100;
    mem[130] = 162'b111111111111111100000000000000000110000000000000001000000000000000001000000000000000000111000000000000000111000000000000001011000000000000000100000000000000000110;
    mem[131] = 162'b000000000000000100000000000000000011000000000000000010000000000000001101111111111111111101111111111111110111000000000000000110000000000000000100000000000000000000;
    mem[132] = 162'b000000000100101011000000000000010000000000000100000101000000000011000111000000000011001110111111111111001101111111111111101110111111111111111110111111111111110111;
    mem[133] = 162'b111111111111111110111111111111111110000000000000000011111111111111110110000000000000000010111111111111111110000000000000110111000000000101000000000000000101111010;
    mem[134] = 162'b000000000000110110111111111111101010111111111111010001000000000000000101111111111111110101111111111111111010111111111111110110111111111111111111111111111111111100;
    mem[135] = 162'b000000000000010000111111111111111110000000000000000001111111111111010110000000000001010110000000000000110111111111111111011110000000000000101011111111111111000100;
    mem[136] = 162'b000000000001100010000000000000110001111111111111101101000000000001000100000000000001000111111111111111000100000000000001010001111111111111000111000000000001010000;
    mem[137] = 162'b000000000000000001111111111111111011000000000000000001111111111111111010000000000000000011000000000000001010000000000100011100000000000110110000000000000101111011;
    mem[138] = 162'b000000000000100000111111111111000110000000000001010011000000000000001011000000000000000001000000000000000011000000000000000110111111111111110110111111111111111000;
    mem[139] = 162'b000000000000011011111111111111100001000000000000000010000000000001000010111111111111110111000000000000110001000000000000010011000000000000111011000000000000011011;
    mem[140] = 162'b111111111111111001000000000000001010000000000000001100000000000000001100000000000000000010000000000000001001000000000000001011000000000000001011000000000000001000;
    mem[141] = 162'b000000000000000101000000000000000001000000000000000100111111111111111101000000000000000010000000000000000001000000000000000000000000000000000100000000000000000000;
    mem[142] = 162'b111111111111111111000000000000000011000000000000000110111111111111111100000000000000000000000000000000000101000000000000000110000000000000000010111111111111111110;
    mem[143] = 162'b111111111111111111000000000000000010000000000000000011000000000000000000111111111111111111111111111111111010111111111111111011111111111111111110000000000000000110;
    mem[144] = 162'b000000000000000111111111111111111101111111111111111001111111111111111000111111111111110111000000000000000110111111111111111001111111111111111100000000000000000110;
    mem[145] = 162'b111111111111111001111111111111111111000000000000000110111111111111111010111111111111111101111111111111111110000000000000000100111111111111111011000000000000001011;
    mem[146] = 162'b111111111111111111000000000000000010000000000000000000000000000000000010000000000000000101111111111111111110000000000000000000111111111111111001111111111111110010;
    mem[147] = 162'b111111111111110110111111111111111001111111111111110011111111111111110111111111111111111010000000000000000000000000000000001001000000000000000000000000000000001111;
    mem[148] = 162'b111111111111110101111111111111111110000000000000000011000000000000000000111111111111111101000000000000000101000000000000001101000000000000001010000000000000000100;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110101111111111111111010111111111111110101;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule