`include "num_data.v"

module w_rom_11 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000000000101000000000110101111000000000000100101111111111011100100000000000001111000111111111110010100111111111100000111000000000000010011000000000001010111;
    mem[1] = 162'b000000000000001010111111100010001111000000000010100101000000000011010010000000000000000001000000001000001000000000000010101100111111010101101110111111110111001011;
    mem[2] = 162'b000000000001001110000000000011011100111111111111110001111111111100110001000000000010010000111111111011011101000000000001001001111111111011011010111111111000000101;
    mem[3] = 162'b111111101100010010111111010101101001111111010011101101111111100100110111111110111010111011111111111101111001111111110110111100111110111111100111111111011000101100;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111110110000110111111111011001011000000000110110010000000000111001000111111111100010101000000000100111010111111111100111010111111110101011011111111110011001010;
    mem[33] = 162'b000000000000101111111111111000111100000000000110110010000000000110001001111111111010100111111111111110101010000000000101111100111111111011110110000000000101000111;
    mem[34] = 162'b000000000001010001111111111101000100111111111010110100000000000011000101111111111110001100000000000000101111111111111100001000111111111111000000111111111110111011;
    mem[35] = 162'b111111110011111101111111111110001001000000000001100111111111111110011000000000000001100110000000000010010001000000000100100101000000000001111011000000001001101101;
    mem[36] = 162'b000000000011100001000000000001000100111111111110101100000000000011010111000000000111110001111111111101010111111111111110110101000000000010110110000000001100101101;
    mem[37] = 162'b000000000000001001111111111111011101000000000000010011111111111101011001111111111010111111111111111110100000111111110110110011111111111111100110000000000001110010;
    mem[38] = 162'b111111111110011011000000000010011011111111111110101110000000001000010011000000000101110111000000000100011100000000000011010000000000000110110000000000000100011101;
    mem[39] = 162'b111111111100100110000000000101111111111111111010101000000000000110000101000000000001001001111111111110011101111111111101011101111111111110011001000000000010111010;
    mem[40] = 162'b000000000110001111111111111110010011000000000000111101111111111100101110111111111110111010000000000100110100111111111110000101000000000110000111111111111101101010;
    mem[41] = 162'b000000000010110000000000000101100011111111111010011000111111111010100101111111111111110101111111111111110011111111111001100000000000000100110010000000000000100011;
    mem[42] = 162'b111111111110001001111111111101000000000000000000001010111111111010101111000000000100010010111111111110000110000000000011011001000000000100010101111111111001110101;
    mem[43] = 162'b000000000110011100000000000011011001111111111111000110000000000111000101000000000011001110000000001010101110000000000001001010000000000001101001111111110111011000;
    mem[44] = 162'b111111111011101010111111111110010110111111111010111101000000000011011010111111111110001110000000000010010101000000001011001110111111111100010000000000001010101010;
    mem[45] = 162'b000000000100101000111111111011000111000000000101011000111111111101011100000000000100111000111111111011001101000000000001011010000000000100110010000000000101010100;
    mem[46] = 162'b000000000110100010111111111011010111111111110101001000111111111101101111000000000100010011111111111111000000000000000001010010000000000011101010111111111001100000;
    mem[47] = 162'b000000001000000111111111111100001010111111111010000010111111111010010110111111111101011001111111111110110010000000000000001111000000000011000000111111110101101111;
    mem[48] = 162'b111111111110000001000000000011010100111111111101001100000000000010101011000000000011000001111111111111110011000000000011000001111111111100010111000000000000010111;
    mem[49] = 162'b111111111011101001000000000000100000111111111000111010111111111001001000111111111101101000000000000010010010111111111011010010111111111110011010000000000000010111;
    mem[50] = 162'b000000000010010010111111111010110101111111110111010011000000000100111110000000000100100111111111111101001010111111111100100100000000000011001000000000000100000001;
    mem[51] = 162'b000000000010000000000000000001010011111111111111100000000000001010110011000000001011010011000000000100111000000000000110110001000000001001011010000000001010010100;
    mem[52] = 162'b000000000111010001000000000110011111000000000001100110000000000010000111000000001000100100000000000101011110000000000111110000000000000111001000111111111110101100;
    mem[53] = 162'b000000001000001011111111111101011010111111111000100011000000000001010000000000000100010110111111111100101110000000000000110010111111111100110011111111111011011100;
    mem[54] = 162'b111111110101000111111111111111111110000000000100101110000000000010100011111111111000101011111111111111111001111111111100010110111111111100011001111111111111101100;
    mem[55] = 162'b111111111001110110111111111101000101111111110111000100111111111100001000000000000001101111000000001010010111000000000000010011000000000000001111111111111111000101;
    mem[56] = 162'b111111111111100101111111110011000100111111111111010100111111111011100011000000000010111111111111111100000010111111111011101001000000000000110101111111111101111100;
    mem[57] = 162'b000000000001100101111111111110001110111111111000000111000000000001001110111111111001110010000000001000101001000000000111000110111111111100111111000000000010010110;
    mem[58] = 162'b111111111001110010000000000110110101000000000010011010000000000100101011111111111111111100000000000000000101000000000011110111000000000001000110111111111100101001;
    mem[59] = 162'b000000001000000111000000000001010110111111111011100011000000000100101110111111111101101000111111111110001010000000000010011101000000000001010110000000000001100010;
    mem[60] = 162'b111111111100101100000000000010010001111111110101101011000000000001111101111111111100010101111111111011111000000000000001001101000000000000100100000000000010010111;
    mem[61] = 162'b000000001000001010111111111100101011111111111000000011111111111111110101000000001001110010111111111001111001000000000010010110111111111111101110111111111011100101;
    mem[62] = 162'b000000000010010110000000000010111001000000000110111010000000000001100111000000000010100111111111111101100011111111111110011100111111111010101000111111111011101001;
    mem[63] = 162'b000000000010101100000000000001111011000000000101011110111111111110010001000000000100110011111111111110101011000000000100001001000000000000010000000000000000101001;
    mem[64] = 162'b000000000011011010000000000011000001111111111110001101000000000011001100111111111110001001000000000000110000000000000101100110000000000110101010000000000000011001;
    mem[65] = 162'b000000000010111000000000000001000101000000000000011001000000000000101010111111110011111111111111111101111110000000000011010101000000001100000011111111111110110000;
    mem[66] = 162'b111111111110100001111111111011100101000000000010011000111111111110101101000000000000111000111111111101011100000000000010001011000000000111111001000000001001100011;
    mem[67] = 162'b000000000000100110000000000011100001111111111100110000111111111101110000000000000000101111000000000110111000111111111111000111111111111101011000000000000100100110;
    mem[68] = 162'b111111111011001100111111111101010011000000000101111011000000000100010101000000000011101000000000000010001100111111111001111001000000000000100100111111110111001100;
    mem[69] = 162'b111111111011111101111111111101011001000000000011100011111111111111000100000000000010001010000000000100110001111111111011000100000000000000000100000000000101101001;
    mem[70] = 162'b000000000101110100000000000011110111000000000010010001000000000010101001000000000000101101000000000101111001111111111001101101000000000001110001111111110111110011;
    mem[71] = 162'b000000000010111011000000000010010011000000000011111100000000000110010000000000000101000111111111111110000110000000000001010011111111111000110011111111111011000011;
    mem[72] = 162'b000000000000110010111111111011000110000000000100010001000000000001001111111111111101111101000000000010111000111111111011101001111111110101001000111111111001101000;
    mem[73] = 162'b111111111001000000111111110011000011111111111000100110111111111110001010000000000011001001000000000001001011111111111110101100000000000100100110000000000010100000;
    mem[74] = 162'b111111111100001000000000000001000001111111111100111111000000000110110111111111111101101110000000000100100011111111111110101101000000000010110100111111111010011010;
    mem[75] = 162'b000000000100000100000000001000000110000000000011110101111111111010100101111111111011001111111111111011100100111111111001001110111111111001110010111111111011110111;
    mem[76] = 162'b000000000101100010000000001000010011000000000011111010111111111110101010000000000100011001000000000101000111111111111110010010000000000001100101111111111101110110;
    mem[77] = 162'b000000000101010101000000000001110010000000000000110100111111111001000100000000000100000011000000000000001000111111111011110010111111111001101010000000000010011111;
    mem[78] = 162'b000000001110101110000000001001110101000000001000100011000000000011010000000000000000110011000000000001110000000000000010111010000000000001001011000000000000111110;
    mem[79] = 162'b000000000001100011111111111011000110111111111011100001111111111101001110111111111111011001111111111110111110000000000010111100111111111111001101000000000001110010;
    mem[80] = 162'b000000000001110000111111111110100111111111111101101100000000000010100010000000000011111011000000000010111010111111111111100110111111111110011000111111111000101111;
    mem[81] = 162'b000000001010110001000000000000111010000000000010110001111111110111010000111111111100011110000000000010000100111111111111001100111111111011000101111111111111001000;
    mem[82] = 162'b000000000010100011111111111000110101000000000111110010111111111110001111111111111101001101111111111111001001000000000101101011111111111011000110111111111011001110;
    mem[83] = 162'b000000000011101010000000000111111100000000000010011010111111111111111101000000000011100101111111111000110000111111111101001011111111111111011011111111111110110100;
    mem[84] = 162'b111111111010010010000000000000101100111111111101110111000000000111001011000000000000100011000000000011000011000000000000100010111111111111000000111111111100100010;
    mem[85] = 162'b000000000111100000000000000000111010000000000010110011000000000001000110111111111100100111111111111010110000000000000010100011111111111101100001000000000100110100;
    mem[86] = 162'b000000000101101101000000000000010101000000000111010101000000000110001010000000001010011001000000001010111100111111111110110101111111111111101010111111111111001110;
    mem[87] = 162'b000000000101110001111111110111011110111111111001101111111111111111110001000000000100001001111111111111011100000000000100010110111111111100110000000000000000011010;
    mem[88] = 162'b000000000001111101000000000100001010111111111101111001000000000000110011000000000000100001000000000101110110111111111111010000111111111010100010111111111001000011;
    mem[89] = 162'b111111111111111011000000000100001011000000000100000101000000000001111111111111111100001101111111111001110100111111111110111000111111111001001100000000000100000110;
    mem[90] = 162'b111111111100011101000000001001100111111111111110001101000000000000100001000000000001011111000000001000110111111111111111101001000000000010000111000000001000010101;
    mem[91] = 162'b000000000001101010111111111111000100111111111100000000000000000011101001111111111110110010000000000110010011111111111001110001000000000010111111000000000010001001;
    mem[92] = 162'b111111111110001010000000000101100001000000000010100000111111111001011000111111111010000100000000000010011011111111111110101100000000000110001011000000000100100011;
    mem[93] = 162'b111111111011100111111111111110000111000000000000101110111111111001001000000000000010100110000000000010010100111111110111101011111111111000001000111111110011000110;
    mem[94] = 162'b000000000001000001111111111101101111111111111100010011111111111110001101000000000010010010000000000110111100111111111111011101000000000010001001000000000001001111;
    mem[95] = 162'b000000000010111111111111111100010101111111111010111010000000000010111010000000000010101101000000000011101111000000000111100010000000000010111100000000000100000000;
    mem[96] = 162'b111111111111111011000000000000001110000000000000010111111111111111110010111111111111111000000000000000000000111111111111101000111111111111111001111111111111110101;
    mem[97] = 162'b000000000000000000111111111111111100000000000000001010111111111111111100111111111111110001111111111111110101111111111111100000111111111111111011111111111111100110;
    mem[98] = 162'b111111111111111010111111111111110111111111111111110110111111111111101010000000000000001111000000000000000010000000000000001010000000000000001011000000000000000000;
    mem[99] = 162'b111111111111101111111111111111110101111111111111110000000000000000001110000000000000000010111111111111111011000000000000001001000000000000001011111111111111111110;
    mem[100] = 162'b000000000000000110111111111111111000111111111111111000111111111111111010111111111111111011111111111111111111000000000000000011000000000000000101000000000000001010;
    mem[101] = 162'b000000000000000011000000000000000001000000000000000110000000000000000001111111111111111110111111111111111111000000000000000000000000000000000011000000000000001011;
    mem[102] = 162'b000000000000010011000000000000010010000000000000000100000000000000000100000000000000000100000000000000001011111111111111111001000000000000001001000000000000001100;
    mem[103] = 162'b111111111111110110000000000000001100111111111111111000111111111111111000000000000000001111000000000000001000000000000000001001000000000000001110000000000000001000;
    mem[104] = 162'b000000000000000100111111111111110100000000000000001001111111111111111100000000000000000110000000000000001100111111111111111100000000000000001100000000000000010001;
    mem[105] = 162'b000000000000000111000000000000000000000000000000000110000000000000000111000000000000000010000000000000000101000000000000000010111111111111111101111111111111111000;
    mem[106] = 162'b000000000000000001111111111111111111000000000000000000111111111111111000111111111111111010111111111111111101111111111111101001111111111111111011111111111111110111;
    mem[107] = 162'b111111111111111000111111111111111010111111111111111100111111111111111011111111111111110011111111111111111011000000000000000101111111111111111110111111111111101111;
    mem[108] = 162'b000000000000001100000000000000001010111111111111111100000000000000000000000000000000001000000000000000000001111111111111101110111111111111111001000000000000000001;
    mem[109] = 162'b000000000000001010000000000000000001000000000000000110000000000000001001000000000000001011000000000000000101000000000000001000000000000000000110111111111111110000;
    mem[110] = 162'b000000000000000010000000000000001010000000000000001010111111111111111001000000000000000111111111111111111101111111111111111111000000000000000000000000000000000101;
    mem[111] = 162'b111111111111111000000000000000000110111111111111111011000000000000000010111111111111111001000000000000001101111111111111111110000000000000000000111111111111111111;
    mem[112] = 162'b000000000000100001111111111111110101000000000000011010000000000000001000000000000000001010000000000000001000000000000000111001111111111111101100000000000000011000;
    mem[113] = 162'b000000000000000111111111111111111101111111111111111110000000000000011001000000000000000000111111111111110000000000000000001100000000000000010111000000000000000000;
    mem[114] = 162'b000000000000010111111111111111111011111111111111111100000000000000000001111111111111111001000000000000000111111111111111111101000000000000001010111111111111111100;
    mem[115] = 162'b000000000000000101111111111111110000111111111111111110111111111111110010000000000000000110111111111111111100111111111111110001111111111111110101111111111111111010;
    mem[116] = 162'b111111111111111110111111111111110111000000000000000101111111111111110100000000000000001010000000000000001111111111111111110110111111111111110000000000000000000010;
    mem[117] = 162'b111111111111111111000000000000001110000000000000000101000000000000001010111111111111111011000000000000000011000000000000001010111111111111111111000000000000000010;
    mem[118] = 162'b000000000000011010000000000000010000111111111111111100111111111111110101000000000000000110111111111111111110000000000000000011000000000000000111000000000000010011;
    mem[119] = 162'b000000000000000100111111111111101011000000000000000000111111111111110011000000000000000000111111111111111010111111111111110100000000000000000101111111111111110101;
    mem[120] = 162'b111111111111111111111111111111111011000000000000010000111111111111111110111111111111110011000000000000000000000000000000001010111111111111111011111111111111110111;
    mem[121] = 162'b111111111111100111111111111111101011111111111111101110111111111111110101111111111111111100111111111111111001000000000000010100111111111111111101000000000000000000;
    mem[122] = 162'b111111111111111011000000000000000000111111111111110010111111111111111110000000000000001000000000000000000011111111111111101010000000000000000110000000000000000000;
    mem[123] = 162'b000000000000000001000000000000001000111111111111111010111111111111111111111111111111111001000000000000000000111111111111111000111111111111110101111111111111111110;
    mem[124] = 162'b111111111111111110111111111111110010000000000000000011111111111111111010000000000000000000000000000000000100000000000000001001000000000000000001000000000000000101;
    mem[125] = 162'b000000000000000010111111111111111010111111111111111100111111111111111000000000000000000111111111111111111101000000000000000110111111111111111100111111111111111110;
    mem[126] = 162'b000000000000000011000000000000001010000000000000000111111111111111111100000000000000001011000000000000001000111111111111101100111111111111110001000000000000000010;
    mem[127] = 162'b111111111111110110000000000000000011000000000000010011111111111111111111000000000000000101000000000000010000000000000000000011000000000000001000111111111111111111;
    mem[128] = 162'b111111111111011001000000000001010010111111111110111001000000000000010110000000000000001101000000000000001110111111111111111101000000000000010101111111111111110111;
    mem[129] = 162'b000000000000000000111111111111110111111111111111111000111111111111111010111111111111110111000000000000000000111111111110111010111111111111101100000000000001100111;
    mem[130] = 162'b000000000000000011000000000000000000000000000000000001000000000000001011000000000000000110111111111111111110111111111111111010111111111111111010111111111111111110;
    mem[131] = 162'b000000000000001000000000000000000000111111111111111000111111111111111001000000000000001000111111111111111111111111111111110111000000000000000010111111111111111101;
    mem[132] = 162'b000000000001100010000000000001000001000000000010110001000000000011100101000000000001110100111111111110101100111111111111110111111111111111100110111111111111111100;
    mem[133] = 162'b000000000000000000111111111111111110000000000000000001000000000000000100000000000000000100000000000000000011000000000010111100000000000010011100000000000011010010;
    mem[134] = 162'b000000000001101011000000000000001101111111111111100101111111111111111111111111111111111110000000000000000011000000000000000000111111111111110111111111111111111111;
    mem[135] = 162'b000000000000100100000000000000010010111111111111001111111111111111111101000000000011101000111111111111001111111111111111110110000000000000010110000000000000101001;
    mem[136] = 162'b000000000001110100000000000000111110000000000010110110111111111111101010111111111111110010000000000000000010000000000000101100111111111111101000111111111111111001;
    mem[137] = 162'b111111111111111110000000000000000100000000000000001100111111111111111101111111111111111011111111111111111010000000000011010111000000000100110101000000000011100000;
    mem[138] = 162'b111111111110110010111111111111111010111111111111010001000000000000000010111111111111111011111111111111111100000000000000000111000000000000001010111111111111111110;
    mem[139] = 162'b000000000000101110000000000000011010000000000000101011111111111110101110111111111111100000111111111110110011000000000000000100000000000001000000000000000001000001;
    mem[140] = 162'b111111111111111100111111111111111010111111111111111111000000000000000011111111111111111001111111111111111011111111111111111010111111111111110001111111111111111111;
    mem[141] = 162'b111111111111111110111111111111111010111111111111111010000000000000000011000000000000000011111111111111111110000000000000000000111111111111111000111111111111111110;
    mem[142] = 162'b000000000000000011000000000000000011000000000000000111111111111111111011111111111111111011000000000000000011111111111111110001111111111111111110000000000000000000;
    mem[143] = 162'b000000000000001011000000000000001000111111111111111111111111111111111011000000000000000101000000000000000101000000000000000011000000000000000110000000000000000000;
    mem[144] = 162'b111111111111111000000000000000001001111111111111111100111111111111111100000000000000000101000000000000000110000000000000000101000000000000000010000000000000000011;
    mem[145] = 162'b111111111111111101111111111111111111111111111111111101000000000000000101000000000000000101000000000000000000000000000000001010000000000000000011111111111111111111;
    mem[146] = 162'b000000000000000101000000000000001000111111111111111101111111111111111100000000000000000001000000000000001011000000000000001111000000000000000001000000000000001001;
    mem[147] = 162'b111111111111111001000000000000001000000000000000000011111111111111111101111111111111111111111111111111111110000000000000000100000000000000001000111111111111111101;
    mem[148] = 162'b111111111111111010111111111111111010000000000000000010000000000000000010111111111111111101000000000000000000000000000000000010000000000000000110000000000000000001;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110111000000000000000000000000000000000000;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule