`include "num_data.v"

module w_rom_6 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000111100000000000000010100100111111111011011010111111111100011010000000000100110011111111111110010110000000000010101001000000000101110101111111110110100011;
    mem[1] = 162'b111111111010000111111111010111111110111111111000001101000000000111111101111111111110110111000000000000011001111111110011000011111111101100011011111111110100000110;
    mem[2] = 162'b111111111110101000000000000001010101111111111100011001000000000010110011111111110111111000111111111010101001111111111110010001111111111011111111111111110010011110;
    mem[3] = 162'b111111100111111000111111100110101011111111111000111001111111010001001011111111010110010100111111101110110001111111011110011101111111100001010011111111101000111110;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111100111100111111110101001110111111110110001101111111111110011101000000000011100001000000000110010000111111110111101101000000000111101010111111110010101011;
    mem[33] = 162'b111111111101010010111111111110111110000000000101110101000000000010010010111111111001111110111111101110101011000000000110101101111111110101010110000000000110001010;
    mem[34] = 162'b111111111000010011000000000000111111000000000010110100111111111100101110000000000111100010111111111110001010000000000011001110000000000100110100000000000001010100;
    mem[35] = 162'b111111111100111011000000000000000111000000000111000000111111111101110110000000000010000010000000000011111111000000000101001011111111111101001101000000000011001100;
    mem[36] = 162'b111111111110000101000000000101001001000000000110011110000000000010110100111111111111010011000000000000110010000000000011110100111111111111001100000000000101101100;
    mem[37] = 162'b111111111111110100111111111100000011000000001100101110111111111101000000111111111111100110111111111010100100111111111111100101000000000001001100111111111100011110;
    mem[38] = 162'b000000000010011101000000000010000101000000000011000000000000000100011001000000001011110101000000000101100010000000000011101001000000000010011011000000000100000110;
    mem[39] = 162'b000000000001011101111111110110101010000000000111110000111111111110110001000000000011000000000000000000100000000000000000011010111111111101101101000000000010011110;
    mem[40] = 162'b000000000111101100000000000001000000000000000100010010000000000001111010000000000011101111000000000100100110111111111001001111000000000011100010000000000010101110;
    mem[41] = 162'b000000000111011101111111111100011001000000000100001010111111111110101101111111111101010110000000001100110001111111111111110111111111111110110011000000000010011110;
    mem[42] = 162'b000000000000000000000000000110111100000000000001111100111111111110001001000000000001000001000000000010011001000000001001011111000000000001000001000000000001101000;
    mem[43] = 162'b111111111110111100000000001000101011000000000100011110000000000111011011000000000010000000111111111011110000111111111010100110000000000010001110111111111000111111;
    mem[44] = 162'b000000001001010111111111111101010101111111111111001110000000000010001101111111111111101111111111111101010111000000000101000010000000000000100111111111111100001000;
    mem[45] = 162'b111111111100010000000000000100111011000000000001010000000000000011000101111111111111100101111111111101000110000000000011110001000000000001000010000000000001011110;
    mem[46] = 162'b111111111110110111000000000000100000111111111110011100000000000111000110111111111000110111000000000001100100111111110100101001111111111100000011000000001010010010;
    mem[47] = 162'b111111111110010000000000001010000101111111110010011001000000000100101100000000000001001111111111111000101101111111111001001111000000000100110101000000000011111000;
    mem[48] = 162'b111111111110110100000000000001010111000000000010011001111111111111110111111111111110101111000000000001111111111111111011111001000000000011001001000000000010111100;
    mem[49] = 162'b111111111110110110111111111111011010000000000001011101111111111110101011111111111100110100111111111001010011000000000010010011111111111100111010111111111111101011;
    mem[50] = 162'b111111111101101000000000000100110110111111111100001111111111111110001111111111111110001101111111111101110010000000000001110010111111110010111111000000000000111110;
    mem[51] = 162'b000000000011001001000000000101010000000000000000100101000000001010101000000000000110100110000000001001000101111111111111101100000000000111101010111111111110111010;
    mem[52] = 162'b000000000101101101000000000000001101000000000000000000111111111111001001000000001001110100000000000011011110000000001000100110000000000100010001000000000001000110;
    mem[53] = 162'b111111111111010101000000000110110110111111111110111000000000000011110001111111111111011010111111110110111001000000000010101011000000000110010011000000000100011001;
    mem[54] = 162'b000000000000100000111111111000000101000000001001110011111111111110100110111111111111010011000000000010001001111111111010101011000000000100001110111111111011101110;
    mem[55] = 162'b111111111101011010000000001011101001111111110010011110111111111110001100000000000101100011000000000001100101000000000010000011000000000010010110111111110011100010;
    mem[56] = 162'b111111111100000111000000000000110010111111111001011100000000000101101110000000000001110001111111111100000101111111110101110111000000000001010110111111111110101100;
    mem[57] = 162'b111111111010011110111111111001101100000000000011001000000000000001000010000000000000100000111111111011100001000000000000111100111111101111001001111111111111101000;
    mem[58] = 162'b000000000101110001111111111110010010111111111110111011111111111001010111000000001000000110111111111010001011111111111110111110000000000101000011111111111111101110;
    mem[59] = 162'b111111111111010001000000000111001001111111111111111000111111110111101111000000000101001110111111110110010011000000000100010110000000000001100001111111111101000110;
    mem[60] = 162'b000000000010011110111111111001111011111111111111000101000000000001011010000000000111010111111111111101000001000000000011110101000000000101111101111111111111001100;
    mem[61] = 162'b000000000001101100111111111110100010111111111011110001000000000100101101000000000010000010111111111000101101000000000011010100111111111001010100111111111011110000;
    mem[62] = 162'b000000000101011111000000000001111110000000000111000110111111111000011100111111111111110000000000000111101111111111111111001010000000000000001111000000000000001000;
    mem[63] = 162'b111111111110101001000000000101000110000000000001000000111111111010001011000000000100010110111111111110101001111111111100001101000000001011000010111111111111100010;
    mem[64] = 162'b111111111110101111000000000010001100111111111101011010000000000001110101000000000000101001111111111100011110111111111010100110111111111100100000000000000000010000;
    mem[65] = 162'b000000000001001001000000000010110100111111111110010010111111111100100101111111111110111101111111111011011010111111111110011011111111111101010110111111111111101100;
    mem[66] = 162'b111111111001110111000000000000101010111111111110110010111111111101000101111111111111001001111111111111100111111111111100100001000000000000110101000000000001111000;
    mem[67] = 162'b000000000010001001111111111110001010000000000010110110111111111110000111111111111111000100111111111101000101111111111110110011111111111110111100111111111110101000;
    mem[68] = 162'b111111111111000111000000000100000101111111111111010101000000000000000000111111111001110000111111111110010111111111111111111000111111111010101011000000000010111010;
    mem[69] = 162'b111111111010001101111111111100001000000000000000011001111111111100111011111111111001010110111111111110101001000000000001100100111111111101100100111111111111001101;
    mem[70] = 162'b111111111110000011111111111101011111111111111111000100111111111101001010000000000000101000000000000100011010111111111000100001111111111010100001111111111001010101;
    mem[71] = 162'b111111111110110010000000000100010101111111111111100010000000000011000110000000000010000100111111111101101011111111111101010101111111111110110010000000000100001101;
    mem[72] = 162'b111111111100101010111111111111001000111111110111011101000000000001101011111111111111001110000000000010011100111111110010010110000000000011100000111111111011101010;
    mem[73] = 162'b111111111001101100111111111111100001111111111101110011000000000000011000000000000011100010111111110110011001000000000001001001000000000001101100111111111001100101;
    mem[74] = 162'b000000000001110110000000000010000010111111111111111010111111111101001100111111111111101100111111111111110011111111111010100110000000000000000001111111111010000101;
    mem[75] = 162'b000000000011001111000000000110011001000000000001001100000000000000100010000000000001110010000000000001101000000000000001100001111111111100010010000000000010101101;
    mem[76] = 162'b000000000100111001000000000011100100000000000011011010000000000110011111000000001001010101000000000111010000000000000010010011000000000011111000000000000000010011;
    mem[77] = 162'b000000000010010000000000000110011010111111111110111111000000000010000011111111111111001110111111111110110000111111111111111010000000000000101100111111111100111100;
    mem[78] = 162'b000000000101101110000000000101001100000000000110100011000000001010001000000000000110010001000000001001010110000000000010100000000000000010101000000000000010101011;
    mem[79] = 162'b000000000000111110000000000101000110000000000000111111000000000011100111000000000000010100111111111101000111000000000101001101111111111100111001000000000101011011;
    mem[80] = 162'b000000000100011111111111111110111110111111111110111000000000000100001010111111111111000100000000000010001100111111111001101001000000000110011101111111111100010010;
    mem[81] = 162'b000000000000100110000000000001110100111111111110101001111111111101100011111111111111001111111111111010011011111111111011101000000000000100001110111111111001010011;
    mem[82] = 162'b111111111101101011000000000000001100111111111110000110000000000100001010111111111100101010000000000001100010111111111000101010000000000101011100111111111000101000;
    mem[83] = 162'b111111111110101001000000000001111001000000000100100001000000000100011011000000000010000011000000000001010100000000000001000001111111111011101010000000000011000010;
    mem[84] = 162'b000000000000111101111111110101010000111111111001000011000000000010100101111111111111100011111111111111110111000000000010010010111111111001010101000000000001010011;
    mem[85] = 162'b111111111110001110000000000000010000000000000001100111111111111110011100000000000011001110000000000010101000000000000000110110111111111111100010111111111100001011;
    mem[86] = 162'b111111111011111101000000000101110101111111111111000111000000000011111000000000000100111010000000000110110111000000000101011100000000001000101000000000000100101101;
    mem[87] = 162'b111111111100111110111111111101100110111111111011000000000000000000011011111111111100101100111111111100011000000000000101100100000000000001111110000000000000100110;
    mem[88] = 162'b111111111111010100111111111010000100111111111100101001000000000010011110111111111110101000000000000100011001111111111010101001111111111110111011111111111110010101;
    mem[89] = 162'b111111111101110001111111111100101110000000000000001011111111111011001001000000000010110100111111111111011100111111111101100110111111111010111110000000000000100100;
    mem[90] = 162'b111111111111001001111111111101101111000000001000010110000000000101001000111111111111101101111111111111110000111111111111101010111111111100011100111111111000110101;
    mem[91] = 162'b000000000001111010000000000000011011111111111100001111000000000001101001000000000110010001000000000010111000000000000011001101000000000100011000000000000001011111;
    mem[92] = 162'b000000000011010010111111111101111100000000000000100010000000000011111101000000000100000101000000000011011101111111111010010100111111110111100100111111111110101111;
    mem[93] = 162'b111111111100000010111111111110001001111111111110011111000000000010010001111111111111111000111111111000100110000000000100011001111111111010011010111111111001111000;
    mem[94] = 162'b000000000001110010111111111111001001111111111111100100111111111010011010111111111001011111111111110111011010000000000011110110111111111011111011000000000101001101;
    mem[95] = 162'b000000000001110111111111111101001100111111111100011110111111111011001010000000000010101011111111111110100111000000000001000110111111111110100110000000000010100001;
    mem[96] = 162'b000000000011000011111111111100010010111111111111001011000000000010110001000000000000001101111111111111011111111111111010111010111111111101100010111111111110010101;
    mem[97] = 162'b111111111101101111111111111110100011000000000010011010000000000000000110111111111111011100111111111110101100111111111110001001111111111101101110111111111110111100;
    mem[98] = 162'b111111111111001010000000000000010011111111111101011101111111111110110000000000000000011011111111111111111001111111111101101110111111111111000110000000000010101011;
    mem[99] = 162'b000000000011000001000000000100111011000000000001100110111111111001000001111111111111011010111111111101111011111111110010010000000000000010100001000000000001100101;
    mem[100] = 162'b000000000000110111000000000000110001000000000010000101000000000100100101000000000001100010000000000011101111000000000010001101111111111111000011000000000001000001;
    mem[101] = 162'b111111111010001100000000000001001001111111111111110110111111111111101110111111111101101110000000000001010001111111111000111101000000000000001001000000000010011100;
    mem[102] = 162'b111111111010100011111111111010010110000000000010110110111111111110100110111111111110001000111111111111100011111111111111110010111111111111011011000000000000010000;
    mem[103] = 162'b111111111100100111000000000000011101111111111001001100000000000010000101000000000000100010000000000001011110111111111111110011111111111100011001000000000001101000;
    mem[104] = 162'b111111111111001000000000000001000011000000000001101101000000000001011011111111111111100001111111111111101111000000000001010011111111111111100001000000000000011100;
    mem[105] = 162'b111111111111101001111111111100011010111111111101111000111111111101110111000000000010111100111111111011000100000000000000011010111111111110010110000000000001001001;
    mem[106] = 162'b111111110111101001111111111001110101111111111001011111000000000010100001111111111100100000111111111100000010111111111010111011000000000010111101111111111101111010;
    mem[107] = 162'b111111111111111001000000000010001001111111111001110010111111111111000000111111111111001110111111111100101101000000000000100001111111111110000101000000000000011110;
    mem[108] = 162'b111111111011000111000000000000111001111111111110111001111111111111001010000000000000011010000000000010011101111111111110010110111111111111001110000000000011111010;
    mem[109] = 162'b111111111110111001111111111011101111000000000001001101111111111100100011111111111101110001111111111111111011111111111110111001111111111111100101111111111100111010;
    mem[110] = 162'b000000000100000010000000000000000010000000000001100111111111111111000111111111111101111001000000000001100001111111111011100011000000000011100110111111111110001100;
    mem[111] = 162'b111111111110011101111111111011110000000000000100001110111111111101010100111111111110101000111111111110110100111111111110010001000000000001000101000000000001100111;
    mem[112] = 162'b000000000101000111000000000010000110000000000111011111000000001111010010000000001000100001000000010011001100000000001110000100000000000100111010000000010000110000;
    mem[113] = 162'b000000000000011001111111111111110010000000000010010110111111111111000001000000000001010011111111111111010000111111111101110010000000000001010001111111111111101001;
    mem[114] = 162'b000000000010110000111111111110011010000000000000010000000000000010001101111111111111100001111111111101000100000000000010101010111111111101110110000000000000111101;
    mem[115] = 162'b111111111111110011000000000000100101000000000001101110111111111110111101111111111110101100111111111110000111000000000001001001111111111110111111000000000010111100;
    mem[116] = 162'b111111111111100100000000000000001001000000000001010101000000000000011000000000000010100001000000000001010000111111111111110110111111111101010000111111111111111101;
    mem[117] = 162'b111111111100100000000000000000011011111111111110100101111111111101100110111111111110010111000000000001001111000000000000101010111111111111110001000000000000001000;
    mem[118] = 162'b111111111010111100000000000010001000111111111100100101111111111110111101111111111111001011111111111111101110111111111010110010000000000001010010111111111110111111;
    mem[119] = 162'b111111111111010011000000000000011011000000000000010100111111111110100101111111111111111100000000000010111001111111111111101110111111111111000000000000000000011000;
    mem[120] = 162'b111111111110101110000000000000100000111111111110110001111111111111011101000000000000001011111111111110001010111111111101100100111111111111111111000000000000010001;
    mem[121] = 162'b000000000011010001000000000010011111000000000011011011000000001100000111000000000110110001000000001100101011000000001010111110000000001000001100000000001111010111;
    mem[122] = 162'b000000000001111000000000000000111011111111111101011000111111111110110011111111111111101010111111111110111111111111111110010011111111111111000000000000000100100110;
    mem[123] = 162'b111111111111110001111111111111000001111111111110100101111111111111111111111111111100010001111111111100010011000000000001101110111111111001111001000000000011000010;
    mem[124] = 162'b000000000010100100111111111101010111111111111010100000111111111110001100000000000000001101111111111111010011111111111111110101000000000010111111111111111111110011;
    mem[125] = 162'b111111111001110011111111111110111010111111111001110010111111111011101101000000000000011110111111111101000110000000000001101011000000000000000101000000000000101000;
    mem[126] = 162'b000000000010001011111111111111110100000000000001100001000000000000000001111111111111010000000000000001110000000000000000011101111111111111000111000000000011011100;
    mem[127] = 162'b111111111111011000000000000000010111111111111101010011111111111111110101000000000000001100000000000001011100000000000001000001111111111101110110111111111111100111;
    mem[128] = 162'b000000000000011000000000000001010100000000000001000010111111111110111011000000000000101101000000000000000110000000000000111011000000000000010111000000000000101000;
    mem[129] = 162'b000000000000000001111111111111111111111111111111111010111111111111111010000000000000000011000000000000000010000000000000001110111111111111001010111111111110111010;
    mem[130] = 162'b000000000000000010111111111111111100111111111111111101000000000000000101000000000000001011111111111111111101111111111111111101111111111111110101000000000000000100;
    mem[131] = 162'b111111111111111110000000000000000101000000000000001010000000000000010000111111111111111011000000000000000011111111111111111111000000000000000110000000000000000001;
    mem[132] = 162'b000000000101000101111111111111000101000000000010100111000000000101000101000000000101010110111111111111110000000000000000001100111111111111110110000000000000001100;
    mem[133] = 162'b111111111111111011000000000000000010000000000000001011000000000000000000111111111111111101000000000000000000000000000000100100000000000010000010000000000101000100;
    mem[134] = 162'b000000000000010110111111111111001111000000000001110010000000000000000111000000000000000000111111111111111010000000000000000011111111111111111111111111111111111101;
    mem[135] = 162'b111111111111111111111111111111110110111111111111100100111111111111000010000000000011111110111111111111100000111111111111000101111111111110100111000000000001111001;
    mem[136] = 162'b000000000000000111000000000000010010000000000001011110000000000001011110111111111111010010111111111111100001111111111111010000000000000010110100111111111111001010;
    mem[137] = 162'b000000000000000011000000000000001011111111111111111100000000000000000101111111111111111001000000000000000010000000000011011011000000000100011000000000000011000110;
    mem[138] = 162'b000000000000101000000000000000100101111111111111011100000000000000000100111111111111111111000000000000000101111111111111111001111111111111111110111111111111110111;
    mem[139] = 162'b000000000000010001111111111111011111000000000000111100111111111111001011111111111111100101111111111111100100111111111111001111111111111111111011000000000011000100;
    mem[140] = 162'b111111111111110100000000000000001001000000000000000100000000000000001011000000000000000000111111111111111110111111111111111110000000000000000100111111111111111001;
    mem[141] = 162'b111111111111111100111111111111111011000000000000001001000000000000000000111111111111111101111111111111111010111111111111110100111111111111110111111111111111111011;
    mem[142] = 162'b000000000000000110111111111111111110111111111111110001111111111111111100111111111111111111000000000000000001111111111111111011000000000000000010111111111111111111;
    mem[143] = 162'b111111111111110100111111111111111110000000000000000100000000000000000101111111111111111011000000000000000000111111111111111101111111111111111100000000000000000000;
    mem[144] = 162'b111111111111110001000000000000001000111111111111111100000000000000000010000000000000001111000000000000000010000000000000000100111111111111111110111111111111111001;
    mem[145] = 162'b111111111111111010111111111111111110000000000000000110000000000000000000000000000000000001111111111111111000111111111111110011000000000000000101000000000000000110;
    mem[146] = 162'b000000000000000000000000000000000010111111111111111001000000000000000110111111111111111000000000000000000011111111111111111101000000000000000000000000000000000000;
    mem[147] = 162'b111111111111111011111111111111110110111111111111111011111111111111110111000000000000001000000000000000000001000000000000000011111111111111111100000000000000001010;
    mem[148] = 162'b111111111111110100000000000000000011111111111111110011111111111111111000111111111111111001000000000000001100000000000000000110000000000000000001111111111111110101;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000001001;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule