`include "num_data.v"

module w_rom_5 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b111111110111100010000000000111011111000000000001011110111111111010001111000000000010100100000000000001101100000000000001011001111111111100110010111111111110000111;
    mem[1] = 162'b111111111110111111000000001001110001000000001000010011111111111100010010000000001001100110111111111110100110111111111011010001000000000001010100000000000001010110;
    mem[2] = 162'b111111111111001111000000000001001101111111111110000011000000000010010011111111111111100101000000000000111010111111111111001010111111111110011101111111111110111011;
    mem[3] = 162'b111111101000010000111111100010010011111111111100000000111111101011111110000000001011010010000000000100100010111111101011010011111111010100100101000000000010100010;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b000000000001110000111111110111000000000000001001001010000000000110111011111111111010011001000000000011010001000000000001100110111111111001010010111111111111111111;
    mem[33] = 162'b000000000000000001111111111110010000000000000001001101000000000011001011111111111110110111000000000010011100000000001000011001111111110011010111000000001000111011;
    mem[34] = 162'b000000000001111101000000000000101011000000000101111010111111111110110000111111111111000000111111111110111110000000000100010010111111111110000101111111111000010000;
    mem[35] = 162'b000000000010110101000000000100111101111111111100110101111111110100110100000000000000011100111111111101110000111111111110110010111111111100000111111111111101100110;
    mem[36] = 162'b000000000100100001000000000110011000000000000001110111111111111110101110000000000000111111000000000110011110111111110110000001000000000001000100111111111101011001;
    mem[37] = 162'b111111111101101000000000000100101101000000000010001001000000000010001010000000000001011111111111111010111000000000000010100111000000000000100100000000000000100000;
    mem[38] = 162'b000000000010010110000000000001011101000000000011010101000000000011000110000000000010000001000000000110010101000000000100010010000000000100000111000000000000011000;
    mem[39] = 162'b000000000110100001000000000010100110111111111000101101000000000000011010111111111111010001000000000100101010111111111100001010000000000011100010111111111000000111;
    mem[40] = 162'b000000000011111010000000001100100001000000000001100011111111111111011110000000000101001100000000000100100111000000000001100011111111111000111001000000000100101001;
    mem[41] = 162'b000000000100101110111111111111100010000000000101101000111111111010110011000000000001100000111111111111101000000000000100000001000000000010101001111111111101100000;
    mem[42] = 162'b000000000001100111000000000001100001000000000000001001000000001000011011111111111101000001111111111111100100111111110111100011111111111110100101111111111111101010;
    mem[43] = 162'b111111111101101100000000000011010000111111111110101110000000000001110000000000000000101000000000000100111100000000000001110001111111111001101011111111111110110101;
    mem[44] = 162'b000000000111010001111111111011111100000000000000010010000000000001011101111111110100111110111111111111111011000000000010100001000000000100101100111111110100110010;
    mem[45] = 162'b000000000010001111000000000000101010000000000100110101111111111010111100000000000000111000000000000100100111111111111110100101111111111110011001000000000000000111;
    mem[46] = 162'b111111111100110110111111111010001111000000000000010000000000000011000111000000000000010111111111111111101100111111111110010111000000000010001011111111111110101111;
    mem[47] = 162'b000000000101011000111111110111101110000000000010011110000000000011011111111111111011110101000000000100101000000000000010001101000000000000111110111111111100110111;
    mem[48] = 162'b000000000010111100000000000010011000111111111010110011111111111110111110111111111101111001000000000100000110111111111101010000000000000010010011111111111011010111;
    mem[49] = 162'b111111110111100001000000000010100000111111111110000000000000000001001111000000000011101010111111110001000111111111111100111110000000001000100101000000000001010111;
    mem[50] = 162'b000000000000101111000000000010001000000000000011101010111111111001010010000000000100000001000000000001001111111111111100001011111111111100011000000000001011000101;
    mem[51] = 162'b000000000010010110000000001000011111000000000101111011000000000100001111000000000010010010000000000011111000111111111111000010000000000010101111111111111100011100;
    mem[52] = 162'b000000000010001001000000001010010011000000000100010110111111111111011000000000000100101100000000000100010110000000000100110001000000000100001001111111111101010001;
    mem[53] = 162'b000000000000001101111111110101111111000000001100111101000000000010101101000000000011101111111111111100010011111111111100001001111111111111011010111111110011010111;
    mem[54] = 162'b000000000001100000111111111100001101000000000110011111111111111100111111000000000000001100000000000110101100000000000011010000111111111010011111000000000011001011;
    mem[55] = 162'b111111111000101000000000000101010010111111111000011010111111111101101010111111111101010001111111111110111101111111111101000000000000000011101100000000000000110110;
    mem[56] = 162'b111111111100101001000000000000010011111111111110000100000000000100011111000000000010111100111111111000110111111111111111011001000000001011010000111111111000101110;
    mem[57] = 162'b000000000011101010111111111011111000000000000011011110000000000010111010111111110101010111000000000110000100000000000001110010111111101110101011000000001000101011;
    mem[58] = 162'b000000000000101010000000000010100101000000000000111101111111111111011111000000000001100101000000000110001000111111111000111101000000000010011010111111111010001010;
    mem[59] = 162'b111111111101100011111111111111001000111111111000011101000000000111010000111111111011101011111111111110011101111111111110101010000000000101011101111111111000101110;
    mem[60] = 162'b000000000010100101000000000001111011111111111001010001111111111011011110111111111110101000111111111111101000000000000000111000000000000001110101111111111100000100;
    mem[61] = 162'b000000000000101110000000000010100111111111111111010101111111111110001010000000000010110111111111111111110100111111111100110101000000000010001001111111111101111010;
    mem[62] = 162'b000000000011110010111111111001100010000000000000001011111111110110111101111111111101100000111111111011011010000000000101000000000000000000000100111111110111111010;
    mem[63] = 162'b111111110111110110111111111111010110000000001010111110000000000000101001000000001010110000000000000001010011000000000100010010111111111111110100000000000011001110;
    mem[64] = 162'b000000000000110110111111111111110110111111111101101111111111111010101110111111111001110001111111111010000100000000000011010111000000000001100111000000000110001010;
    mem[65] = 162'b111111110111101110000000000001001001000000000000101001111111111111011000000000000001100110111111111110111100111111111111100010000000000011011011000000000000111110;
    mem[66] = 162'b111111111011100101111111111110110100111111111110110111000000000010001110111111111000111001111111111100010011111111111011100101111111111100100011000000000110111010;
    mem[67] = 162'b000000000100001000000000000001100101111111111110111100000000000000110100000000000010101100111111111111101010000000000001100001000000000000011010111111111101110110;
    mem[68] = 162'b000000000000110110111111111011001000111111111100011000000000000000000110000000000010110010111111111111010001111111110100010110111111111011001101111111111111100100;
    mem[69] = 162'b111111111111000011000000000000010100000000000001001010111111111011001000111111111010011110000000000011111100000000000011011101111111111001111100000000000001111101;
    mem[70] = 162'b000000000011011001000000000001110011111111111100010011111111111111011001111111111111100110111111111011111101000000000001111110000000000100011000000000000011000110;
    mem[71] = 162'b111111111111010101111111111010010001111111111110101011000000000011001111000000000001110011000000000001000001111111111100010010111111111101101101111111111100010000;
    mem[72] = 162'b000000000111111011111111111111010011000000000010111011111111111100011010000000000010011000000000000100010110000000000000000101000000000001100011111111111110100101;
    mem[73] = 162'b000000000000010000000000000000111000000000000000101011111111111111000010111111111100001100111111111111101111000000000001111011111111111110110001111111111101000101;
    mem[74] = 162'b000000000100000110111111111011100001111111111010011101111111111000000100000000000010100111111111110101001000111111111111111110111111111110100011111111111000111010;
    mem[75] = 162'b111111111101111110000000000000000011111111111111001110000000000001001100000000000000010100111111111111100101111111111110100011000000000000100100111111111110101000;
    mem[76] = 162'b111111111110101101111111111111110110111111111110101011000000000010001010000000001001011011000000000110110111000000000010000010000000000101111111000000000010111011;
    mem[77] = 162'b000000000000111111000000000001100110111111111100001100000000000011111010111111111110110000000000000011110111111111111010001011000000000001010111111111111000100000;
    mem[78] = 162'b000000000101000101000000000100111000000000000010110011000000000101111100000000001001111001000000000110000010111111111111110010000000000010111001000000000011100010;
    mem[79] = 162'b000000000000111001000000000011010001111111111101111101111111111101110010111111111101000000000000000100111110111111111111100011111111111111000111111111111101000000;
    mem[80] = 162'b000000000001101011111111111110100000000000000001000001000000000010001110000000000010010001111111111111011101000000000001111101111111111111000100111111111110101010;
    mem[81] = 162'b111111111011011011111111111111001101111111111111111011000000000000001010000000000011100010000000000000001011111111111001100111111111111111100001000000000001001000;
    mem[82] = 162'b000000000001101000111111111110011000111111111100000110111111111100111000111111111111110001000000000000010101000000000110000011000000000011111010000000000100100100;
    mem[83] = 162'b000000000111111011111111111101110010000000000100011111000000000001011011111111111111011100111111111101000101000000000111011010111111111110110001000000000111010101;
    mem[84] = 162'b000000000001111000000000000010011001111111111010010010111111111110101111111111111000101111000000000001001001000000000001111000111111110111101011111111111101001000;
    mem[85] = 162'b111111111111010011111111111100101111000000000001001011000000000100111110000000000001000111111111111110001101111111111101010111111111111111011100111111111001000101;
    mem[86] = 162'b000000000001000110000000000100100001000000000000111111000000000110101000000000000110000010000000000110000101000000000001010011000000000110100100000000000110100010;
    mem[87] = 162'b111111111111010110111111111111100010111111111110111110111111111101001111000000000010110100111111111011101111000000000000111111111111111111110001000000000001111100;
    mem[88] = 162'b111111111111011011111111111100100000000000000010010101111111111011111101111111111101000011111111111111111000000000000010011101111111111111010101000000000100000010;
    mem[89] = 162'b111111111101100101000000000000100100000000000001010110000000000010111011111111111110110000000000000010000000111111111110110000111111111100011010111111111100000111;
    mem[90] = 162'b111111111101001101000000000000101110111111111110010110111111111011111010111111111101101010000000000001011011000000000000111001111111111110011110000000000011011101;
    mem[91] = 162'b111111111110101001000000000100011100000000000000010111111111110110101100000000000000001000000000000110110100000000000101000010000000000111001101000000000111110110;
    mem[92] = 162'b111111111101111100000000000001000000000000000011111100000000000011110100000000000010101100000000000000110010111111111010101101111111110110111000111111111111010111;
    mem[93] = 162'b111111111111111011000000000010111010111111111100101011111111111101111110000000000010100000000000000000110101000000000101010110111111111101010001111111111000111000;
    mem[94] = 162'b000000000010010001000000000000100101111111111010101101111111111100001111000000000011010101111111111101010010111111111111101001000000000011100001111111111101111011;
    mem[95] = 162'b000000000111010110000000000000100100000000000110011100111111111111100101000000000011010010111111111111011000111111111101111100111111111111101000111111111110101001;
    mem[96] = 162'b111111111110101001111111111110010010111111111010101101111111111101100111111111111110001101111111111100110101111111111100100101111111111111011110000000000001101111;
    mem[97] = 162'b111111111110110111000000000000011011111111111100100011000000000001001010111111111100101010111111111111011010111111111111100101000000000000101010111111111110110111;
    mem[98] = 162'b111111111111111111111111111110111101111111111110001011000000000001010001111111111100110100111111111101011100111111111111100011000000000000011100000000000011110001;
    mem[99] = 162'b000000000000111100111111111100000110000000000001110001111111111111100011111111111101111010111111111000001101000000000000101100111111111011110000111111111111011101;
    mem[100] = 162'b000000000000111111000000000011101000000000000010110100111111111110110110111111111111111111111111111101101011111111111110010011111111111110011001000000000000011100;
    mem[101] = 162'b000000000010101110000000000000010000000000000000101101111111111101001011111111111110000011111111111100111001111111111100111000111111111110001010000000000000000000;
    mem[102] = 162'b111111111110100000111111111111001110000000000000101101000000000001001010000000000000110011000000000000111101000000000011110001000000000001011111000000000100001011;
    mem[103] = 162'b111111111110100111111111111100111100000000000010011001111111111100001000111111111101110110111111111110100110111111111101110011000000000001100110000000000011111001;
    mem[104] = 162'b111111111110100000111111111110101000000000000010100111000000000001000100000000000001000111000000000001110101111111111101011001000000000001001011000000000010101101;
    mem[105] = 162'b111111111011011101000000000001010000111111111101101000111111111101011110111111111111111111000000000000010010111111111111100001111111111100000111111111111111011111;
    mem[106] = 162'b111111111111010111111111111101011111111111111011000111111111111101110110111111111111001011111111111001000011000000000001101011111111111100110100000000000100001111;
    mem[107] = 162'b000000000000110000000000000000000101111111111000110010111111111111000010111111111110111100111111111110011011111111111100011000111111111111111010111111111111000101;
    mem[108] = 162'b111111111100001001111111111111100000111111111101011111000000000001111101000000000000110011111111111110011001111111111001100110000000000010111011111111111110101111;
    mem[109] = 162'b111111111100110001000000000000110001111111111111011101111111111111001010111111111101111111111111111111100000000000000000100000111111111101001011111111111101000101;
    mem[110] = 162'b111111111110101101111111111101111100111111111101000001000000000000011011000000000000001000000000000001100100111111111010001011111111111110110111000000000010100000;
    mem[111] = 162'b111111111101100101111111111110000011000000000000010110111111111111111010000000000000110001000000000001100101000000000001110110111111111011011100111111111111010110;
    mem[112] = 162'b000000000011000001000000001010100010000000001001010000000000000111101111000000001010000010000000001000100011000000000010110111000000001001011110000000001011101001;
    mem[113] = 162'b111111111000101101111111111011010001111111111101010001000000000001011000000000000001101000000000000000100011000000000000101000111111111110110001000000000010010101;
    mem[114] = 162'b000000000000011001000000000000011110000000000010001111111111111011101011000000000000110101111111111111000001000000000000110011000000000000000100111111111011000101;
    mem[115] = 162'b000000000011011001000000000000111110111111111100100011111111111110111110111111111111110001111111111101100111111111111111010111000000000001011000111111111110010101;
    mem[116] = 162'b111111111110100111111111111101101011111111111100111010111111111111100110111111111101110111000000000010000010000000000000001010000000000000111001111111111111000000;
    mem[117] = 162'b000000000001101111111111111111111000111111111110101010000000000001010100000000000001010111000000000011001000111111111100011110000000000000110111000000000000111001;
    mem[118] = 162'b111111111101010100111111111110100011000000000000110100000000000000100111111111111111011110111111111110000101111111111110000011111111111110011101000000000001100001;
    mem[119] = 162'b111111111001110100111111111111000100000000000000011100111111111110010110111111111111011111000000000011001110000000000001001100000000000000101010111111111111111000;
    mem[120] = 162'b000000000010111101000000000001100111000000000011001101111111111100110110111111111101100010111111111100100011000000000001001100111111111110101110000000000000111010;
    mem[121] = 162'b000000000100001111000000000110010110000000000110100110000000001010101000000000001010101001000000000111101001000000000011110111000000001101001011000000001010101100;
    mem[122] = 162'b111111111110010011000000000000010010000000000000100001111111111111110101111111111110001110000000000010100111111111111111101111111111111101110011111111111111111000;
    mem[123] = 162'b000000000001001011111111111110111110111111111101111001111111111111101101000000000000011010111111111110010110111111111111001000111111111001110001000000000001001001;
    mem[124] = 162'b111111111111000011111111111111100101111111111110010101111111111011001001111111111100001001000000000001100001000000000001010101000000000000100010111111111100111110;
    mem[125] = 162'b111111110101010000000000000000110011111111111100010001000000000001100000111111111110100110000000000000100000111111111100011010000000000001111111111111111111010000;
    mem[126] = 162'b000000000000011111111111111110001010111111111110000101000000000000110110111111111111111101111111111111110110000000000000000011000000000001011110111111111101110101;
    mem[127] = 162'b111111111111011111111111111111001010111111111110100101000000000001101110000000000000011101111111111101111100111111111101101111000000000000110010000000000000001000;
    mem[128] = 162'b111111111111011000111111111111011110000000000000111111111111111111111011000000000000010110111111111111011111111111111111100010000000000000010011000000000000011110;
    mem[129] = 162'b000000000000000001111111111111110100111111111111110101000000000000001000111111111111111011000000000000000000111111111111010100111111111111010111000000000010000101;
    mem[130] = 162'b000000000000000001111111111111111110000000000000000010000000000000001010111111111111111101111111111111110111111111111111111101111111111111111000111111111111111000;
    mem[131] = 162'b111111111111111101111111111111111001111111111111111011000000000000000000000000000000001001000000000000000100000000000000010010000000000000001001111111111111110100;
    mem[132] = 162'b000000000100010111111111111111110100000000000010100110000000000100110000000000000011010100000000000000001100000000000000110001111111111111101101111111111111110011;
    mem[133] = 162'b000000000000000110000000000000001100000000000000000010111111111111111101000000000000000001000000000000000111111111111111101010000000000011011101000000000100110010;
    mem[134] = 162'b111111111110010100111111111111001100111111111111111011000000000000001101111111111111110000000000000000010100111111111111111000000000000000000110000000000000000100;
    mem[135] = 162'b111111111111000110000000000000011001000000000000000100000000000000011011000000000010110010111111111111111000111111111111111000000000000000011100000000000000010100;
    mem[136] = 162'b111111111111101000000000000001100111000000000001011001000000000000001111000000000001010100000000000000010000000000000000100101000000000001011100000000000000110100;
    mem[137] = 162'b000000000000000010111111111111111010111111111111110101111111111111110000111111111111111000000000000000000000000000000100000000000000000011010100000000000101001110;
    mem[138] = 162'b000000000000001001000000000000010000111111111111111001000000000000000100111111111111111101111111111111111000111111111111111000111111111111111100111111111111101110;
    mem[139] = 162'b111111111111011011111111111111011000000000000010001001111111111111011011111111111111010100000000000000010111000000000000000100111111111111100110000000000000000001;
    mem[140] = 162'b111111111111110000000000000000000001111111111111111010111111111111110110111111111111110011000000000000000111111111111111111011111111111111111010111111111111111011;
    mem[141] = 162'b111111111111111010000000000000000101111111111111110111111111111111110101111111111111111111000000000000000001111111111111110001111111111111101011111111111111101111;
    mem[142] = 162'b111111111111111111000000000000000000000000000000000000111111111111111000111111111111101011111111111111110011000000000000001010111111111111111100111111111111111000;
    mem[143] = 162'b000000000000000001111111111111111011111111111111111010111111111111110111111111111111111111000000000000000001000000000000000001111111111111111011000000000000000100;
    mem[144] = 162'b111111111111111101000000000000000000000000000000000100000000000000001000111111111111110111111111111111111000111111111111111001000000000000000001000000000000000010;
    mem[145] = 162'b000000000000010001000000000000011001000000000000010010000000000000000000000000000000000000000000000000011010000000000000000010111111111111110001111111111111111011;
    mem[146] = 162'b000000000000000000000000000000000001000000000000000110000000000000001001111111111111111011000000000000000000000000000000010000000000000000001000000000000000000000;
    mem[147] = 162'b111111111111100101111111111111111100111111111111111110111111111111111001000000000000001101111111111111111101000000000000010011000000000000000110000000000000001101;
    mem[148] = 162'b000000000000010000000000000000001011000000000000000010000000000000000010000000000000000000000000000000011110000000000000000011000000000000001011000000000000001010;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111101000000000000000110000000000000001000;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule