`include "num_data.v"

module w_rom_23 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000100100001000000000000001011000000000110010100000000000001111011000000000110010110111111111111110100000000000001101000000000000000001001000000000100010111;
    mem[1] = 162'b111111011001110010111111011100110001000000000001010110111111111100010110000000000001110111111111110101111001111111011110101101111111001110010011111111111011110011;
    mem[2] = 162'b000000000010101011111111111100111110000000000001011001111111111111000101000000000010000100000000000000010101111111111000001100000000000001101001111111111101010101;
    mem[3] = 162'b111111111000011000111111111100010100000000000001000110111111110100011101111111100011111101111111110100000110111111101001001001111111011111000101111111101010100110;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111110101010001000000000110101101111111111100000001000000000000111100000000000011110100111111111110111001111111110111000010111111110110011001111111111100111110;
    mem[33] = 162'b000000000011110101000000000100101000000000000111010000111111111111111101000000000101101101111111111110110100111111111010111010111111111000111100111111111100000111;
    mem[34] = 162'b000000000011110001000000000110000011000000000001001100000000000001001100111111111101001101111111111011001110111111111001001111111111111100110111000000000111000001;
    mem[35] = 162'b111111111101111001111111111111110100111111111010000011000000000110010011111111111110001111000000000110111100111111111011001110111111111100010110000000000010010100;
    mem[36] = 162'b000000000101011101111111111101110000000000001000001111000000000010001011000000000000011110111111111110100101000000000111110101111111111101010000000000000100110101;
    mem[37] = 162'b111111111101101101000000000010101000000000000010111011000000000100011011111111111110111101111111111101001000000000000001101011111111111110010100111111111101001000;
    mem[38] = 162'b000000001000000010000000000001111011000000000011011110000000000010110000000000000001110110000000001010110111000000000100101101000000000100001001111111111101100110;
    mem[39] = 162'b111111111111001000000000000100010111111111111100101011111111111110011001000000000000001101000000000100000001111111111110101110111111111011100000111111111101000111;
    mem[40] = 162'b000000000000111100000000000111000100000000000010011111000000000010010110111111111101100001000000000001010101000000000011111100111111111011000101000000000011110101;
    mem[41] = 162'b111111111011000000111111111000110000000000000011100100000000000110011000111111110101011111000000001001101101000000000000110011111111111100100000111111111010101000;
    mem[42] = 162'b000000001001001010000000000000111100000000001010000100111111111100010010111111111100010010000000000101011000111111111101001011000000000000110000000000000010111100;
    mem[43] = 162'b000000001001001110000000000011010010111111111101100010000000010000100110000000000001011111000000000100000100000000000011011011000000000010001111111111111010000011;
    mem[44] = 162'b111111111100111010000000000100000111111111111001010110111111111111001100000000000001111000111111111111101000000000000100010010111111111100101010111111111110000011;
    mem[45] = 162'b111111111111101010000000000001001110111111111011101111111111110100100101000000000000101100111111111011111001111111111010011110000000000010011011111111111001101010;
    mem[46] = 162'b000000001010100000000000000010110000111111110111111111111111110110001111111111111111110011111111111110011001000000000100010001111111111011101010111111110110110010;
    mem[47] = 162'b000000000111100100000000000000011111111111111101110101111111110111010001111111111011111110111111111111110001000000000100011100000000000100010000111111111111100010;
    mem[48] = 162'b111111111110010000111111110011010000111111111110010111111111111110010011000000000011011100000000000101011101111111110101110001111111111111110110000000000001100001;
    mem[49] = 162'b000000000101001011111111111111000110111111111011000101000000000001111001111111111001011101111111111000011000000000001000001111000000000010101100111111111100000011;
    mem[50] = 162'b000000001010111000000000000111000011111111111011000101111111111001101011111111111111100101111111111110111001000000000101100011111111111011111011111111111001110111;
    mem[51] = 162'b000000000010100111000000000101100001000000000110001010000000000011001100111111111111101001000000000111011011111111111110100010000000000001001010000000000111010011;
    mem[52] = 162'b000000000001101001000000000101001000000000000110111001000000000110010110000000000010011110000000000001101101111111111011001111111111111100010101000000000001100011;
    mem[53] = 162'b000000000100110011000000001000111010111111111001100111111111111110010010111111111101111011000000000100000100111111111110001101111111111011010110000000000000010001;
    mem[54] = 162'b111111111110010011111111111101110011111111111001011001111111111101000101000000000101111101111111111111111010000000000011100011111111111110001001000000000001000111;
    mem[55] = 162'b000000000011011001000000000100001011111111111101011111111111111111001010111111111101101100000000000001111111111111111100001111111111111101110111000000000111100100;
    mem[56] = 162'b111111111100100110000000000011010110111111110111011010111111111111001000111111110111101000000000001000111011111111111010011001000000000011011011111111111111001001;
    mem[57] = 162'b000000000001010001000000000011101010000000000010111110000000000010100001000000000011111000111111111111010100111111111010110011111111111111010111111111111111001011;
    mem[58] = 162'b000000000100010000111111111110111010000000000110000100111111111110111001000000000101111011000000000101101100111111111100010001000000000000001111000000000010101110;
    mem[59] = 162'b000000000010001110000000000001110101111111111001110110111111111101100011111111111101100011000000000111100110111111111111101011000000000101001010000000000000001000;
    mem[60] = 162'b000000000001110011000000000000010101000000000000100111000000000110110010111111111111001111111111111000111110000000000001110111000000001000000011111111111101101000;
    mem[61] = 162'b000000000001110000000000000101001110000000000111010010111111111100011111111111111101001010111111111110111011111111111110011011111111111101000011111111110101101011;
    mem[62] = 162'b111111111011100100111111111011101000111111111010110110000000000111010001111111111111010010111111111110110001000000000110010110000000000001101000111111111100100111;
    mem[63] = 162'b000000000001000111111111111100101101111111111101010001000000000001100000000000000010000100000000000010110101000000000101101100000000000010011110000000000100110010;
    mem[64] = 162'b111111111111000010000000000010000010000000000100000001111111111100101111000000000011100101111111111110101000111111111110011010000000000010000100000000000000011100;
    mem[65] = 162'b111111111101111110111111111111111010111111111000111111111111111001111101111111111011000011000000000000100100000000000100000101000000000101000111000000000001100101;
    mem[66] = 162'b000000000001010000000000000010101111111111111100101100000000000000100111111111111011100110111111111111010110000000000101001100111111111100100110000000000001101011;
    mem[67] = 162'b000000000100000010111111111111000011000000000100110001111111111001000011111111111100111100000000000000010001111111111110100110000000000001101101000000000010111001;
    mem[68] = 162'b111111110111001111000000000000000000000000000111001001111111111010000000000000000010001100111111111100110101111111111010111000000000000000000111111111111101001110;
    mem[69] = 162'b111111111001101101111111111111000111111111111111111011111111111001101100000000000000001011000000000001010011000000000011010110000000000111000010000000000000100000;
    mem[70] = 162'b000000000000111011111111111100110001000000000111011000000000000110101011000000000000101100111111111110000100000000000001001001000000000001111110111111111011101010;
    mem[71] = 162'b000000000000011000111111111101100001000000000000111111111111111111100000111111111111111011111111111111101000000000000011010001111111111011001100111111111100101010;
    mem[72] = 162'b111111111111110110111111111110000011000000000011101001111111111111011101111111111010011011111111111011111001111111111101101111111111111111100100111111111111011001;
    mem[73] = 162'b000000000000110100111111111101000111000000000000101000000000000010010110111111111110011000111111111111010100000000000101101010000000000010001010111111111100001001;
    mem[74] = 162'b111111111101011011000000000000110010111111111110100101000000000010000001111111111110010001111111111001011000111111111100101110000000001000000011111111111101110101;
    mem[75] = 162'b000000000000110000000000000011100111000000000100001000000000000000111101000000000010010011111111111111100110111111111101110111000000000011010110111111111000011111;
    mem[76] = 162'b000000000100010011000000000111001101000000000010110111000000000100000100000000000101101001111111111111010011000000000110100011000000000111000001000000000110011110;
    mem[77] = 162'b000000001000110001000000001000010100111111111101001101111111111110110011111111111011110111000000000001000100111111111000000001111111111001100011111111111111110100;
    mem[78] = 162'b000000000101110100000000000101010001000000000101111001000000001010001100111111111110011001111111111011110101000000000101100101000000000110001100000000000001001001;
    mem[79] = 162'b000000000010000110111111111111100000111111111010101111000000000001100111000000000101101100111111111110100110000000000000001000111111111111110110000000000010101001;
    mem[80] = 162'b111111111010001000000000000111110110000000000110000000111111111101011010111111111110000000111111111001101010000000000000011010000000000010011100000000000011010111;
    mem[81] = 162'b000000000001100001111111110111111101111111111111011000111111111011110110111111111100010001111111111110000111000000000000101110111111111001011101111111111111100010;
    mem[82] = 162'b000000000001011110111111111011110001000000000001111100111111111110110010111111111100000101000000000101011111000000000010001110000000000000111110000000000011110110;
    mem[83] = 162'b111111111110010110000000000100011110000000000000011101111111111010111111000000001000011110111111111101001011000000000100001010000000000011011001111111111111101101;
    mem[84] = 162'b000000000100110101111111111010011000111111111011000100000000000001001101111111111100101101111111111101001010000000000011001000111111111100011001111111111111001100;
    mem[85] = 162'b111111111110111100111111111110010100111111111100101000111111111110101011111111111011010011000000000011101000000000000011111011111111111111101110111111111111100001;
    mem[86] = 162'b000000000011011110000000000111011011000000000110010110000000000110011100000000000011001111000000000001010011000000001110100111000000001100111011000000000111111000;
    mem[87] = 162'b111111111101101101000000000011000000111111111101000001000000000100100011000000000010010100000000000001000010111111111011010100000000000000101110111111111111011010;
    mem[88] = 162'b000000000001000000000000000001011000111111111110110000000000000000010011111111111101010000111111111110001001111111111001011000000000000000111100111111111010001100;
    mem[89] = 162'b111111111010111111000000000000110010111111111101000011111111111111100111111111111110101000000000000100010011111111111111110110111111111100011110111111111110011111;
    mem[90] = 162'b111111111101011100000000000010110001000000000101111101111111111001110111111111111111111100000000000001110110111111111101110001000000000010011111111111111011001100;
    mem[91] = 162'b111111110101100110000000000000101011000000000101001101000000000100011111000000000000110001000000000010100010000000000101010111000000001000011110000000000001110110;
    mem[92] = 162'b000000000100111000111111111111011000111111111110101100000000000001010000000000000000011100111111111100110001000000000011100011111111111000111100111111111111000001;
    mem[93] = 162'b000000000000100111111111111001000011111111111100101110111111111111011001000000000000001100111111111110100001000000000010100001111111111110000010000000000101000101;
    mem[94] = 162'b111111111010011010111111111110101011000000000010011000000000000000011111111111111111010011111111111011011011000000000000100101111111111011010000111111111101011101;
    mem[95] = 162'b111111111101101001000000000001000011111111110110100010111111111111001111111111111101001101111111111111100101000000000100110111000000000110001111000000000000001000;
    mem[96] = 162'b000000000000000100000000000000001111111111111111111101111111111111100011000000000000011110000000000000011001000000000000000100000000000000000001111111111111111010;
    mem[97] = 162'b111111111111110001000000000000000101000000000000010010000000000000010010111111111111111101111111111111110101111111111111100000111111111111110111000000000000001111;
    mem[98] = 162'b000000000000010101000000000000000100000000000000101010111111111111111101000000000000011101111111111111111001000000000000000101000000000000001000000000000000000111;
    mem[99] = 162'b111111111111111010000000000000001101000000000000011110111111111111101001111111111111110111000000000000001011111111111111110110111111111111110011111111111111110100;
    mem[100] = 162'b000000000000100010000000000000001011000000000000000111000000000000010001000000000000001111000000000000000100000000000000001100000000000000001010000000000000000100;
    mem[101] = 162'b111111111111100001111111111111110001000000000000010010000000000000001001000000000000010000111111111111110000000000000000001000000000000000000011000000000000011110;
    mem[102] = 162'b000000000000000100111111111111110100111111111111101101000000000000010100000000000000010000000000000000010011000000000000010010000000000000010001111111111111111110;
    mem[103] = 162'b000000000000010011111111111111111001111111111111111000000000000000011100000000000000000110000000000000000001000000000000000101000000000000000101111111111111110101;
    mem[104] = 162'b000000000000000011000000000000001010000000000000011111000000000000000111000000000000001001000000000000000001111111111111111111111111111111101101111111111111111011;
    mem[105] = 162'b000000000000001101000000000000011001000000000000011010111111111111111011000000000000010001111111111111111000000000000000010101000000000000000111111111111111101101;
    mem[106] = 162'b000000000000000101000000000000010000000000000000001110000000000000000011000000000000010000000000000000001010111111111111111101000000000000011001000000000000001000;
    mem[107] = 162'b111111111111110100111111111111110000000000000000000001000000000000001011000000000000000011000000000000000101000000000000010010000000000000010000000000000000000111;
    mem[108] = 162'b000000000000001010000000000000011100111111111111101111111111111111110001000000000000010011000000000000010000000000000000000010000000000000001010000000000000000101;
    mem[109] = 162'b111111111111111100000000000000000001000000000000001000111111111111110100000000000000000100111111111111110011000000000000010101111111111111111011000000000000000110;
    mem[110] = 162'b000000000000010010000000000000000001000000000000001010000000000000010100111111111111111100000000000000000111111111111111111111000000000000000010000000000000001101;
    mem[111] = 162'b111111111111011011111111111111101110111111111111111111111111111111111011111111111111111111000000000000010000000000000000000110000000000000010111000000000000000000;
    mem[112] = 162'b000000000000101111000000000000001010000000000000111000000000000000001110000000000000010010000000000000011010111111111111100110000000000000010010000000000000101000;
    mem[113] = 162'b000000000000010100111111111111101001000000000000001000000000000000011001000000000000011000000000000000011101111111111111111001111111111111111010111111111111111100;
    mem[114] = 162'b000000000000010100111111111111110010111111111111101101000000000000000111000000000000001101000000000000000110111111111111110010111111111111110010111111111111111100;
    mem[115] = 162'b111111111111101001000000000000000100111111111111111101000000000000000000000000000000011111000000000000100001000000000000000111111111111111110111111111111111101111;
    mem[116] = 162'b111111111111100100111111111111111110000000000000000111111111111111010010000000000000000110000000000000011111111111111111101011111111111111101110111111111111100110;
    mem[117] = 162'b000000000000000001000000000000010111111111111111101010000000000000000110000000000000010001000000000000100011000000000000001100000000000000010100111111111111101001;
    mem[118] = 162'b000000000000101010000000000000010111111111111111111111000000000000011000000000000000001110000000000000000101000000000000000100000000000000010010111111111111110011;
    mem[119] = 162'b111111111111111110000000000000001000000000000000011000000000000000001011000000000000000011000000000000010001000000000000001100000000000000010111000000000000001110;
    mem[120] = 162'b000000000000000111000000000000001010000000000000010100000000000000000111000000000000001010000000000000101110000000000000010111000000000000001001111111111111111011;
    mem[121] = 162'b111111111111111111000000000000000100000000000000100001000000000000000000000000000000001011000000000000000101000000000001110100000000000000001010000000000000011111;
    mem[122] = 162'b111111111111110100111111111111011011111111111111111001000000000000001110000000000000001010111111111111111011111111111111011111111111111111110000000000000000000010;
    mem[123] = 162'b000000000000011000000000000000000011000000000000001011000000000000010101000000000000000101000000000000000010000000000000001001111111111111110110111111111111111101;
    mem[124] = 162'b000000000000000110000000000000001010000000000000000010000000000000001010111111111111111110000000000000000000000000000000000101000000000000010000000000000000000100;
    mem[125] = 162'b111111111111111010111111111111101111111111111111110010000000000000001000000000000000001101111111111111110011000000000000001010000000000000001010111111111111111110;
    mem[126] = 162'b000000000000101000111111111111110101000000000000010011000000000000000001000000000000001011000000000000010000000000000000010000000000000000000010111111111111101011;
    mem[127] = 162'b111111111111111011000000000000001001111111111111110000111111111111100010111111111111111111111111111111101110111111111111110110111111111111111011111111111111100101;
    mem[128] = 162'b000000000010011001000000000100111010000000000100111011000000000101011000111111111111101101111111111111101010000000000000000110111111111111111101111111111111111011;
    mem[129] = 162'b000000000000000010111111111111111011000000000000000001000000000000000010000000000000000100111111111111111110000000000000001001111111111111011010000000000000010011;
    mem[130] = 162'b000000000000000010000000000000001010111111111111111110111111111111111011111111111111110111000000000000000100111111111111111110000000000000000011000000000000000100;
    mem[131] = 162'b111111111111111010000000000000000011000000000000000011111111111111111000111111111111111110111111111111111001000000000000000111000000000000000100111111111111111011;
    mem[132] = 162'b000000000000110111000000000000011111000000000000011110000000000000000011000000000000000001111111111111111001111111111111101010111111111111100110111111111111111000;
    mem[133] = 162'b000000000000000100000000000000001000111111111111111101000000000000001010000000000000001110111111111111111101111111111111011110000000000011101010111111111111011100;
    mem[134] = 162'b000000000101011010000000000100111000000000000100100011000000000000001100111111111111111101000000000000001001111111111111110110000000000000000110111111111111111110;
    mem[135] = 162'b000000000000001010000000000000100000000000000001000010111111111111111011000000000000000010111111111111110010000000000001111010111111111111010100000000000011000101;
    mem[136] = 162'b111111111111110101000000000000000001000000000000000100000000000000001000000000000000000101000000000000000001000000000000001101000000000000000110000000000000000110;
    mem[137] = 162'b111111111111111010000000000000001100111111111111111111000000000000000001000000000000000010111111111111111001111111111111111110000000000000000101000000000000000010;
    mem[138] = 162'b000000000000000000000000000000000100111111111111111111000000000000001001000000000000000010000000000000000110000000000000001001000000000000000011111111111111111010;
    mem[139] = 162'b111111111111111100000000000000000000000000000000001101000000000000000100111111111111111010000000000000000010111111111111111110111111111111111011111111111111111100;
    mem[140] = 162'b000000000001111101000000000011000010000000000010011001000000000000000100111111111111110110111111111111110010000000000001010001111111111111110011111111111100001101;
    mem[141] = 162'b000000000000000010111111111111111110000000000000000000111111111111111111111111111111111110111111111111111001000000000011011111000000000100111011111111111111111010;
    mem[142] = 162'b000000000011000001000000000011010110000000000011100111111111111111111011111111111111111111111111111111111001111111111111111000111111111111111111000000000000000010;
    mem[143] = 162'b111111111111110010000000000000010110000000000000001110000000000000101110111111111111011001000000000000100001111111111111111010000000000000001010000000000011110011;
    mem[144] = 162'b000000000000000000000000000000000001000000000000000010111111111111111000111111111111111100111111111111111011000000000000000011111111111111110010111111111111111110;
    mem[145] = 162'b111111111111111100111111111111111111000000000000000100000000000000001011111111111111111001111111111111111111000000000000000000000000000000000001000000000000001000;
    mem[146] = 162'b111111111111111101000000000000000010000000000000000101000000000000000001000000000000000010000000000000000001111111111111111010000000000000000011000000000000000000;
    mem[147] = 162'b000000000000000011000000000000001011000000000000000010000000000000000001111111111111111110111111111111111100000000000000000000111111111111111101111111111111111100;
    mem[148] = 162'b000000000000000101111111111111110101111111111111111111000000000000000101111111111111111101000000000000000001000000000000000110000000000000000011000000000000000001;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110111111111111111100000000000000001000;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule