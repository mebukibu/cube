`include "num_data.v"

module w_rom_0 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000110100000000000000010110011111111111010111011000000001100101100111111111110101100111111111000110110000000000000110010000000000001110000111111111101000111;
    mem[1] = 162'b111111101111100101111111111010110001111111110110110110111111110110111101000000000111011001000000000000101100111111111101111110111111111010001001111111111011000000;
    mem[2] = 162'b000000000000001010000000000010001110111111111111111101111111110111011011111111111011001000000000000000011010000000000010100011000000000111111101000000000101000101;
    mem[3] = 162'b000000000101111100000000000100110101000000000000000111111111100111000111000000001010101110111111101010110110000000001000110000000000000010100101111111111111101000;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111110010001111111111111111010111111111000101110000000000000101000000000000000010101111111111000000100000000000001001001000000000100110010111111111111110111;
    mem[33] = 162'b111111111100101001111111111100100010000000000100110010111111111100000110111111111111101000000000000100000011111111110110110011111111111001000011000000000110100010;
    mem[34] = 162'b111111111011010100111111111111010110111111111100010111000000000011011000111111111011001110111111111010110010111111111001000111000000000111100110000000001010100110;
    mem[35] = 162'b111111111000000111111111111011111000111111111001101110111111110111010111111111111100110111000000000110111110111111111100111110111111111111100101000000000100010001;
    mem[36] = 162'b111111111111101010000000000010110001000000000010111110000000000100110111111111111101101101000000000101011100111111111000001000000000000011011000000000000101111001;
    mem[37] = 162'b000000000100011011111111111100000010000000000100000000000000000000101101111111111100011001111111111010111110111111111000011111000000000010111000000000000000001100;
    mem[38] = 162'b000000000101110101000000000001110011111111111111101011000000000000100110000000000101011000000000000010110100000000001000000001000000000001100110000000000011001110;
    mem[39] = 162'b111111111110010010111111111100100110111111110011100000111111111011110001000000000011000101111111111111100010000000000000101011111111111111111100000000000010011101;
    mem[40] = 162'b000000000001010011000000000000100001000000000011000010111111111101001001000000000101011111000000000001110010000000000101001010111111111100100010111111111011000100;
    mem[41] = 162'b111111111101101101111111110110000100111111111101000001111111111101011100000000000100011011111111111111111101000000000100010000111111111111010110111111111110000100;
    mem[42] = 162'b111111111011001111000000000000011001000000000010011110000000000010000011000000000010011110000000000100010000000000000010100011111111111110010100111111111101000000;
    mem[43] = 162'b000000000100101100111111111111001010000000000000000000111111111101100100111111111011100001000000000100001110111111111111110100000000000110010000000000000001110100;
    mem[44] = 162'b000000000100000011111111111111100010111111111010000001111111111101011100111111111110011000000000000010101101000000000001100101111111111010000000111111111101100000;
    mem[45] = 162'b111111111111011011000000000000010101000000000101101111000000000011010100000000000010101000000000000000000010111111111110010011000000000001100111111111111000100110;
    mem[46] = 162'b000000000010001111000000000110111101111111111101001000111111111000000101111111111101111100000000000101111111111111111111011001111111111010111011111111111110101100;
    mem[47] = 162'b000000000001111010000000000001100100111111111000000011000000000011110001111111111100101100000000001000101000000000000101011000000000000000010000111111111010000111;
    mem[48] = 162'b111111101110111001000000000001010100000000000010111011000000000111010011111111110111101100000000000100110010000000000010111101000000000001001011111111110110111110;
    mem[49] = 162'b111111111010001100111111111111010111000000000011010000000000000100010100111111111110101111111111111110000011111111110010001010111111110110110010111111111100000001;
    mem[50] = 162'b111111111100101110000000000100010010111111111111001011111111111111000101111111111100110001111111111100110001000000000001110010000000000011001100111111111010101011;
    mem[51] = 162'b000000000011000100000000000011101001000000000000001100000000001000000100000000001111010000000000001010000000000000000100010111000000001011111111000000001010001110;
    mem[52] = 162'b111111111110000011000000000001011101111111111110001110000000000110111010000000000101000100000000000101110000000000000110001011000000000100000000000000000101001010;
    mem[53] = 162'b111111110110111010000000000010011100111111111010101011000000000001110100111111111010110101000000000011110100000000000000101110000000000000110000000000000111001011;
    mem[54] = 162'b111111110100100101111111111110100010000000000100111111000000000010001001111111111101100100000000000000010000000000000100100101000000000110001000111111111000010101;
    mem[55] = 162'b000000001001101010000000000000100010111111111001011100000000000010011100111111110011110101111111110110101111111111111010010001000000000100101101111111111100110110;
    mem[56] = 162'b111111111000001010000000000011000001000000000001101011111111111000001111111111111101000100000000000101100110111111111100110110000000000011111110111111111001111010;
    mem[57] = 162'b000000000001110001111111111100010011000000000000101110000000000011110101111111111111010001111111111110011011111111111110111011111111111100110000000000000001111110;
    mem[58] = 162'b000000001000111010111111111111001001111111111101101100000000000011110101111111111001110101111111110111100010111111111101101111111111111110010100000000000111100111;
    mem[59] = 162'b111111111000101100111111111010101001000000000110000101000000000101011000111111111011001000111111111000100011111111110111000010000000000000111110111111111100001101;
    mem[60] = 162'b111111111100000100000000000000100000111111111111001100000000000010111000111111110110100010000000000000010000000000000010100101111111111010100011000000000110100110;
    mem[61] = 162'b000000000010011001111111110111100000111111111111001011000000000000010010111111111110101010000000000010000101111111111100010001111111110111100001000000000010100110;
    mem[62] = 162'b000000001000010111111111111111001011111111111010101110000000000001110010000000000111010010111111111010111001111111110101010111111111111000010011000000000100001011;
    mem[63] = 162'b000000000010001111000000000011111011000000000010100111000000000100100011111111111100001110000000000000001100111111111101110000111111111100111101000000000011000100;
    mem[64] = 162'b111111111100001101111111111011100010000000000010000100000000000011100011000000000011011010000000000100101110000000000001100010111111111101100101111111111110100110;
    mem[65] = 162'b000000000110101000111111111010101110111111111111100101111111111010100100000000000000101000111111111110100011000000001001110001000000000001011011000000000111001000;
    mem[66] = 162'b000000000001011010000000000101110111000000001000100000000000000010010100111111111101100010111111111011111100111111111110011000111111111010000011000000000000010000;
    mem[67] = 162'b000000000000101000111111111100000001111111111101110101111111111101111001111111111101101110111111111110111001000000000110011011111111111110010010111111111101111110;
    mem[68] = 162'b000000000000101011111111111101111111000000000001001111000000000011110110111111111111001101111111111011100101111111111101100000111111111110100100111111110111010101;
    mem[69] = 162'b000000000100000011111111111010001010000000000001001111000000000011111000111111111011001110000000000110110000000000000010110011111111111110001101000000000000101101;
    mem[70] = 162'b000000000000011100000000000101101000111111111111101010000000000010111110000000000100000010000000000001101001111111111001111100111111111110000001111111111011111100;
    mem[71] = 162'b000000001000101101000000000100111010000000000000110010000000000110001110000000000100111011111111110101001110111111111100100101000000000010011001000000000101100001;
    mem[72] = 162'b111111111010001010000000000001001011111111111010001010000000000000000100111111111011010000111111111101111111111111111110000010111111111011101000000000000000001101;
    mem[73] = 162'b111111111001010111111111111011010100111111111110011001111111111101111011111111111011111111111111111100001011111111111010111110111111111111010000111111111111000100;
    mem[74] = 162'b111111111111001000111111111110000010111111111010100101000000000100100110111111111001110111111111111101010000000000000100110000111111111100010010111111111011100001;
    mem[75] = 162'b000000000001011011000000000110100011000000001010100011000000000100001011111111111100110110111111111110110111111111111111011001000000000000010011000000000000000100;
    mem[76] = 162'b000000000100111010000000000001100001000000000111100101111111111110000110111111111110111111000000001000001011000000000001010011000000000010000011000000000111010010;
    mem[77] = 162'b000000000001111100000000000010100110000000000010001101111111111110110101000000000000100101000000000000110101111111111111100111111111111010111011000000000000110110;
    mem[78] = 162'b000000000111110100000000001000011001000000000111011110000000000011111001111111111111101011000000001000001010000000000001000110000000000011010000000000000101111101;
    mem[79] = 162'b111111111001011100000000000110011101000000000001111010000000000000101101000000000110110101111111111110001000000000000000101001111111111111011111000000000110000000;
    mem[80] = 162'b111111111110101110000000000110101111111111110101011001000000000000101010000000000100100010111111111011101110000000000011010111111111111110101000111111111100100000;
    mem[81] = 162'b000000000000011100111111111010000110000000000010110001000000000000000110000000000001101010000000000101000010000000000001111111111111111000110111111111111110010001;
    mem[82] = 162'b000000000111100110000000000010111101111111111100000001000000000001110000111111111111101101000000000010000100111111111100011100000000000000010100000000000100111111;
    mem[83] = 162'b000000000001001101000000000101101110000000001000100101111111111111011100000000000110101010111111111111111110000000000010001011000000000100101001000000000100001100;
    mem[84] = 162'b111111111110000100000000000001000110111111111111100110000000000010110011111111111100010010111111111110101101000000000100000010000000000001000100111111111010101010;
    mem[85] = 162'b000000000000001100000000000001011111000000000110101110111111111101111110111111111010010001000000000011100111000000000001000101111111111111110100000000001000000101;
    mem[86] = 162'b111111111110011000111111111110010100000000001001100001000000001000001011000000001001000000000000000111111110000000000001011101000000000001010100000000000101100111;
    mem[87] = 162'b000000000011001010000000000000101000000000000010101000000000000010110001111111110111010100111111111100101000000000000010010001111111111110101100111111111100110010;
    mem[88] = 162'b111111111011111001111111111110010001000000000100000010000000000010100110111111110100101011111111111011100010111111111101011011000000000000101001000000000000101000;
    mem[89] = 162'b000000000001000011111111111110000000111111111110111110000000000100011011111111111110000110111111111001001010111111111011001100000000000111110011000000000001010100;
    mem[90] = 162'b000000000110111010111111111111100100000000000000000101111111111010110001111111111101011011000000000011000100111111111110000010000000000011000001000000000000100100;
    mem[91] = 162'b111111111111010001111111111000000100111111111010101001000000000111111001000000000110000011000000001001111001000000000010100011000000000001100001111111111111011000;
    mem[92] = 162'b000000000011001100111111111010111100111111111110101011111111111000011000111111111111001111000000000110010110111111111011010011000000000100100011111111111100110010;
    mem[93] = 162'b000000000001110000111111111011110011111111110110011001000000000011101100111111111011001101111111111100011110000000000110110010111111111011101101000000000001101110;
    mem[94] = 162'b000000000000000011000000000001001000111111111100111110000000000010110011000000000000011110111111111011101001111111111011000010000000000000001110000000000100110000;
    mem[95] = 162'b000000000000111111111111111100110010111111111110100100111111111110010011111111111011010011111111111111110001111111110101000101000000000000000100000000000010111001;
    mem[96] = 162'b000000000010000110111111111011011110111111111011100101111111111110110010111111111111001101111111111111100000000000000010110010111111111110100111111111111111111110;
    mem[97] = 162'b111111111101010101111111111111110010111111111110011000111111111111111001000000000000110011111111111011001101000000000000001111111111111111001000111111111100100011;
    mem[98] = 162'b000000000001000011111111111101001001111111111111010110111111111111100111111111111111000010000000000000101000111111111110110000111111111110100111111111111110110001;
    mem[99] = 162'b111111111111011001000000000000111011000000000101000001111111111101111010111111111110000010111111111101011101000000000010000110111111111100010001111111111111100001;
    mem[100] = 162'b111111111101111111000000000011110001000000000010110011000000000011001101000000000000000111000000000001111011000000000011000101111111111100011010111111111110010101;
    mem[101] = 162'b000000000000100111111111111110100011111111111011110100000000000000010000000000000000010000111111111110010110111111111100001010000000000001000000111111111110100101;
    mem[102] = 162'b111111111101010100000000000001000111111111111111110011000000000000001011000000000100000111111111111101111011000000000001010111000000000000010110111111111101001101;
    mem[103] = 162'b111111111101011110111111111111000110000000000011100111111111111111100111111111111111110101111111111101011001000000000001101111111111111100101010111111111110001111;
    mem[104] = 162'b000000000000011010000000000001010110111111111111110111000000000010011111111111111101110111111111111111011110000000000000001010111111111101000111111111111110111100;
    mem[105] = 162'b111111111101110100111111111110010111111111111110101010000000000000011011111111111111100001000000000000100101111111111111000001111111111111011100000000000000000010;
    mem[106] = 162'b111111111110000100111111111110011000000000000000110011111111111101100001111111111101000011000000000000011111000000000000001111111111111111001110000000000001011100;
    mem[107] = 162'b111111110111011110111111101110110100000000000010100111111111110111110000111111111000001110111111111101111011111111111110001100111111111001101011111111111110100001;
    mem[108] = 162'b111111111110110010111111111111000110111111111111010110111111111101010001111111111111001011111111111111100010111111111110100011111111111111100001000000000001011001;
    mem[109] = 162'b111111111110110101000000000001101110111111111110110111111111111111100110000000000010100101111111111011111101000000000000001011111111111111101011111111111110000001;
    mem[110] = 162'b111111111101001111111111111110111000000000000100011011111111111101000011000000000001000110000000000001010010111111111111001100111111111101110001111111111111010101;
    mem[111] = 162'b000000000001110001000000000000010111000000000001010010000000000000000110111111111101010100000000000001110111000000000001101010000000000000011001000000000000001101;
    mem[112] = 162'b000000001000101101000000001000010000000000000101011100000000001011110111000000001001001010000000001000110111000000001001001101000000000101001111000000000111101000;
    mem[113] = 162'b000000000000101001000000000001000101111111111100001101111111111110100000111111111111110010000000000000001111000000000000001000111111111110101111111111111101111000;
    mem[114] = 162'b000000000000010111000000000001101000000000000010011100111111111110110010000000000000000010111111111110101000111111111111011000000000000000001001111111111111010101;
    mem[115] = 162'b111111111011000100111111111111000010111111111111001001111111111111110111000000000000101000000000000010001000000000000000011000111111111101011000111111111010100001;
    mem[116] = 162'b111111111111110101000000000010110011000000000000101110000000000000000011111111111111001111111111111111101011000000000000001011000000000010000001111111111101101011;
    mem[117] = 162'b111111111100101111000000000000011000111111111110111101000000000000111100111111111111101100111111111111000011000000000000110101111111111001100000000000000000100001;
    mem[118] = 162'b111111111111000100111111111111101110111111111101100010111111111111100000111111111101111101000000000001001010111111111111101011111111111111101111111111111110000000;
    mem[119] = 162'b000000000011010001111111111111001001111111111111110110111111111110101101000000000000101111111111111110011001000000000001011001000000000000010001000000000001111111;
    mem[120] = 162'b111111111111101101111111111110101011111111111101100001000000000000000110000000000000010011111111111101011110111111111101111100111111111101000001000000000000001000;
    mem[121] = 162'b000000000100111110000000000101001001000000000000111001000000001001100110000000000111111110000000000100101110000000000110011110000000000110011000000000000011000000;
    mem[122] = 162'b111111111101101101000000000000000110111111111101110010000000000000000111111111111111011100111111111110101000111111111111110101000000000000100100111111111110000011;
    mem[123] = 162'b000000000011010101111111111111001110111111111100001100000000000000010100000000000000100100111111111111000001111111111100000100000000000001100011111111111111011000;
    mem[124] = 162'b000000000001010100000000000000010000000000000001000001000000000000011010111111111101101011000000000000101010111111111101010001000000000010000010111111111000111110;
    mem[125] = 162'b000000000010111111000000000000110101111111111110110000111111111110011110000000000001000011111111111011001100111111111111110000111111111011110011111111111100111010;
    mem[126] = 162'b000000000000100111000000000000011001000000000000111011111111111101111110000000000000110011111111111111111000111111111111010000111111111111010010000000000001000010;
    mem[127] = 162'b000000000000000011111111111110010100000000000000101001111111111111001010111111111111011111111111111111100101000000000000000110111111111110100011000000000000000011;
    mem[128] = 162'b000000000000100101000000000000010111000000000000010010000000000000011010111111111110110001111111111111110001000000000000000011000000000000010110111111111111010010;
    mem[129] = 162'b111111111111111100000000000000000000111111111111110101111111111111110111111111111111111100111111111111110001111111111111010110111111111110100101111111111110101110;
    mem[130] = 162'b111111111111111000000000000000000110000000000000000100000000000000001010000000000000000111000000000000000010000000000000001101000000000000000011111111111111111000;
    mem[131] = 162'b111111111111111100000000000000001001111111111111111110000000000000000001111111111111110111111111111111110011111111111111110000111111111111110000111111111111110001;
    mem[132] = 162'b000000000011111110000000000000101010000000000000100011000000000011011000000000000001111001000000000001100110111111111111010001000000000000000011111111111110111100;
    mem[133] = 162'b000000000000000100111111111111111111000000000000000111000000000000001001000000000000010101000000000000000111111111111111110110000000000011010101000000000100000110;
    mem[134] = 162'b000000000000100000111111111111010110111111111111011010000000000000000111000000000000000001111111111111111000111111111111111011000000000000000001000000000000000011;
    mem[135] = 162'b111111111111110001111111111111010001111111111111100111000000000000010010000000000010101011111111111111100100000000000000001110000000000001100010111111111111101110;
    mem[136] = 162'b000000000011010111111111111110000101000000000010011010111111111111110000000000000000111010111111111111111110000000000000111010000000000000101100111111111111001111;
    mem[137] = 162'b111111111111110100111111111111111110111111111111110110000000000000000110111111111111111111000000000000001010000000000010010111000000000010001101000000000100010101;
    mem[138] = 162'b111111111111110000000000000001101011000000000001010001000000000000001001000000000000001000111111111111111101111111111111110000000000000000000010111111111111111011;
    mem[139] = 162'b000000000000011111111111111111100011000000000000011100111111111110111111111111111111011010111111111111111001111111111111101001000000000001011111000000000011010110;
    mem[140] = 162'b111111111111111000000000000000001000000000000000001000111111111111111111000000000000000101111111111111111011111111111111111110111111111111111010111111111111110000;
    mem[141] = 162'b111111111111111011111111111111111011000000000000010001000000000000000011111111111111111111111111111111111110111111111111110100111111111111111101111111111111111010;
    mem[142] = 162'b111111111111111110000000000000000111000000000000001111111111111111110111111111111111111111111111111111111011000000000000000001000000000000000010111111111111111010;
    mem[143] = 162'b000000000000000110111111111111111111000000000000000000000000000000000000111111111111111001111111111111111000111111111111111101111111111111110111111111111111111111;
    mem[144] = 162'b000000000000001010111111111111110100111111111111110110111111111111111010111111111111110000111111111111111010000000000000000000000000000000000101000000000000010001;
    mem[145] = 162'b111111111111111110000000000000000110000000000000001101000000000000000110000000000000001111111111111111111110000000000000001111000000000000000110000000000000000000;
    mem[146] = 162'b000000000000001010000000000000001101000000000000001001111111111111110111111111111111111111000000000000010000111111111111111011000000000000000111000000000000000000;
    mem[147] = 162'b111111111111110010111111111111111111111111111111111000111111111111111100000000000000000010000000000000000110000000000000000001000000000000000010000000000000001100;
    mem[148] = 162'b111111111111111101000000000000000000000000000000000000000000000000001000000000000000001010000000000000010001000000000000001100000000000000001110000000000000010001;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111111111111111110;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule