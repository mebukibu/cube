`include "num_data.v"

module w_rom_12 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000000111110111111111100100100000000000001010011000000000001000001111111111101110101000000000110101010000000000011111001000000000101100111111111110000111011;
    mem[1] = 162'b000000000010000101111111111001001111111111010110010001111111111001010100111111111001000101000000000010111110000000000011111010000000001101010100111111001001110110;
    mem[2] = 162'b111111111011110100111111111111011100000000000001011101000000000000010001000000000011100001111111111011000000000000000001000101111111111111111001111111111100010011;
    mem[3] = 162'b000000001110110110000000000011010110111111111000111100000000000100110101000000000000010110111111110101101100000000000011010100000000000000101001111111101101111011;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b000000001001110010111111111110101000111111111111101110111111111101001101000000000001110011000000000010010011111111110011011001111111111010110100111111111101101011;
    mem[33] = 162'b000000000011000111111111111010101001000000000001110001000000000010111100111111111111001110000000000111010010111111110011010011000000000001100111000000000001101001;
    mem[34] = 162'b111111111011111011111111111110011000111111111110010011111111111001111110111111111110000110000000000110011110111111110111010010111111110101000011111111111101110001;
    mem[35] = 162'b000000001000000000111111111110100111000000000101001000111111111001110010111111111001010000000000000111010001111111111101010100000000000011010101111111111100011100;
    mem[36] = 162'b000000000100101100000000000010000011000000000101001011000000000100010101000000000101110001000000000110110000111111111101011011000000000000100101111111111111101110;
    mem[37] = 162'b000000000011000110111111111111010000111111111001001001000000000100011001111111111100011010000000000000101110000000000110100111111111111111010100111111111101111101;
    mem[38] = 162'b000000000111111000000000001010010111000000000011010000000000000111001010000000001001001000000000000110110000000000000010001001000000000001110111111111111111110100;
    mem[39] = 162'b000000000110110000000000000101101100000000001000000010000000000100000101000000000000110001111111111110010010111111110101000011000000000001011100000000000011001100;
    mem[40] = 162'b000000000111010011000000000110100000000000001010101010000000000010111110000000001011000010000000000100011001000000000101010011000000000101111111000000000000110011;
    mem[41] = 162'b000000001010101100000000000000101011000000000000111000000000001010001100000000000110110010111111111111001100000000000110100001000000001001000001000000001000110010;
    mem[42] = 162'b111111111100010000000000000110111000000000000110001010000000000000100011000000000001111001000000000011000111111111111110000111111111110111110001000000000100111100;
    mem[43] = 162'b111111111111100111000000000001010000000000000010001011000000000011111111000000000001100010000000000110000000111111110111010110000000000011110011111111111101111000;
    mem[44] = 162'b111111111011000011000000001001110110000000000010011101111111111101100101111111111100110100000000000100110101111111111010100111111111111110010100000000000010001001;
    mem[45] = 162'b000000001001110001000000000001010000000000000011010101111111111000110011000000000010000000000000000001110000111111111111011001111111111011100010111111111110101011;
    mem[46] = 162'b000000000001000110000000000110101011000000000101110101111111111110100100000000000100011110111111111101010111111111110101010011000000000000000011000000000101001110;
    mem[47] = 162'b111111111000101100000000000111101010000000000101010100111111111110010000111111111110010000000000000100011101000000000000011010111111111010010110111111111101011110;
    mem[48] = 162'b000000000111000001000000000011111111111111111110111010111111111101000111111111111101011001111111111111111011000000000010000000111111111001110100000000000000011100;
    mem[49] = 162'b111111111111100101111111111010001110111111111100101110111111111110101010111111111110100000111111111001001111000000000101011011000000000000110011000000000010011000;
    mem[50] = 162'b000000000011001101000000000010001111000000000010101100111111111010011100000000000000100011111111111111011111000000000111001110111111111100101111000000000010111110;
    mem[51] = 162'b000000001111001010000000001111001101000000001010001111000000001011001110000000001011100011000000001011111011000000000111110011000000000101101001000000000011010000;
    mem[52] = 162'b000000001001010111000000001001000111000000000110011100000000000101101101000000001000001000000000000111010001000000000010010011000000000101111010111111111101000110;
    mem[53] = 162'b000000000001111001111111111100110101000000000101001010111111111110100000111111111110100001000000000101100111111111111001110101000000000001100110111111111110001101;
    mem[54] = 162'b000000000010111000000000000101001001111111111111011101111111111101011011000000000010000110000000000000101010111111111101111101000000000110001101111111111011000000;
    mem[55] = 162'b000000000111011101000000000011000010000000000101100100111111111001110100111111110111010111111111111100110101000000000110000101000000001000010110111111111110000101;
    mem[56] = 162'b000000000110011101111111111110100100000000000011110011111111111011111011000000000010000001111111111010111001111111111000100010000000000110010101111111111011111110;
    mem[57] = 162'b000000000110100010111111111001111110111111111011111111111111111011010101111111111011110110000000000011111001000000000011011001111111111010010111000000000100000010;
    mem[58] = 162'b000000000110111000000000000011010101000000000011001001000000000000011111000000000010110100000000000011100101000000000000110100000000000100001111111111111110110100;
    mem[59] = 162'b000000000010001010000000000001001011000000000000101011000000000000110100111111111001011010111111111110011100000000001001000101111111111100011101111111111001000110;
    mem[60] = 162'b000000000010110101000000000011010010000000000000100011111111110101101111111111111101101110000000000100110100111111111011101000111111111111110111111111111110111001;
    mem[61] = 162'b000000001010110110111111111101010101111111110100001100000000000000001000000000000100001011111111111100011101000000000010111000111111111111001111000000001010001100;
    mem[62] = 162'b000000001001101011000000000111101000000000000011000101111111111100011111111111111010011110000000000000110001111111111011111110111111111000110011111111110111100000;
    mem[63] = 162'b000000001000101010000000001100111101000000000101000001000000000000000100000000000011000111000000000100010100111111111110100101000000000101101011111111111101101101;
    mem[64] = 162'b000000000011111111000000000000001001111111111101110100111111110111101100000000000110000111000000000000100101000000000110100000111111111011100101111111111101010010;
    mem[65] = 162'b000000000000011110000000000101001000111111111000000011000000000010101111111111111111100100111111111111011001111111111111011001111111111001101011000000000001110100;
    mem[66] = 162'b000000000000001000111111110110011110111111111101000010111111111100000100111111110110111010000000000000110010111111111011101100000000000001100000111111111010001000;
    mem[67] = 162'b111111111100001010000000000100101010111111111011010111000000000011011011111111111111011001111111111101000000000000000001011100000000000000111111000000000000101100;
    mem[68] = 162'b000000000010000110111111111110011111111111111110111111111111111011000011111111111101001000000000000000111010111111111011110011111111111110000011000000000101011011;
    mem[69] = 162'b111111111110000111000000000010101000000000001000011011111111111101110110111111111100011101000000000001000100000000000000010100000000000010011110111111111111100010;
    mem[70] = 162'b000000000000100000111111111101111101000000000010111101111111111010010101111111111111001110000000000011110111000000000011001010111111111101111001111111111100111101;
    mem[71] = 162'b000000000011000011000000000000110001111111111101110110111111111100100101111111111110000101111111111100101101000000000010101101000000000001011101111111111101001101;
    mem[72] = 162'b000000000011010110000000000000000000111111111101111111000000000010100100111111111110100011000000000001001101111111111000000110111111111110110001111111111101000001;
    mem[73] = 162'b111111111110100111000000000001011100111111111011011100000000000001011000000000000000100110111111111110011011111111111111111001000000000010000101111111111110010000;
    mem[74] = 162'b111111111110100000111111111011100101111111111011000001111111111100100100000000000011101000111111111101011110111111110111011101000000000100011001111111110111110011;
    mem[75] = 162'b111111111110110000111111111111101011000000000001011000000000000011001101000000000001011101111111111110110011000000000000010000000000000001010101111111111111010000;
    mem[76] = 162'b111111111111111111000000000010010011111111111111001111000000000010010110000000000011100101000000000011100001000000000001100111000000000110110100111111111110110100;
    mem[77] = 162'b000000000100110011111111111111001010111111111111000111000000000001000000111111111110100010111111111101111010111111111000101001111111111110010111000000000000111101;
    mem[78] = 162'b000000001000100001000000000001111001111111111110110000000000000100011010000000000101111111000000000101111111000000000100111000000000000001000100000000000101100011;
    mem[79] = 162'b000000000101100001000000000000111110111111111100011011111111111110001010000000000000010000000000000010001100000000000110000001111111111101000110111111111101001000;
    mem[80] = 162'b111111111110100000000000000001001111000000000011000111000000000101101111111111111011111101111111110111100001000000000100011001000000000001110100111111111111001010;
    mem[81] = 162'b111111111110101100000000000011011001000000000001101101000000000000110100000000000000001101111111111101001100000000000001010101000000000000011100000000000000110111;
    mem[82] = 162'b000000000010010100000000000000000111000000000100001100000000000111100001000000000110011111000000000101101000000000000010000000111111111001011101000000000001000011;
    mem[83] = 162'b000000000011101110000000000001100010000000000011011101000000000101100011111111111110110110000000000100000111000000000001100100000000000000000101111111111101000110;
    mem[84] = 162'b000000000011101011111111111110011111000000000110001111000000000010010010111111111101101010000000000011110010000000000010110010111111111011100001111111111001011010;
    mem[85] = 162'b000000000101011101111111111111011001111111111100000100000000000100011111111111111111011011111111111111001011000000000110000000000000000000110100111111111100101100;
    mem[86] = 162'b000000000011000000000000000001100100000000000010010010000000000111010100000000000100000111000000000011111001000000001000111111000000000001111101000000000011011011;
    mem[87] = 162'b111111111011110010000000000000001011111111111101101111000000000010001010111111111110011010111111111011101011000000000010100011111111111110011101111111111110111101;
    mem[88] = 162'b000000000010011000000000000101000001000000000101010111111111111101111111111111111111011100111111111111011110000000000010110110111111111100011010111111111111011010;
    mem[89] = 162'b111111111101001100111111111101011111111111111111111000000000000010001010111111111111000001000000000001100111111111111111010101111111111111000010111111111111100111;
    mem[90] = 162'b000000000000100011000000000100001000000000000001010000000000000010100110000000000001010010000000000001000011000000000011011001000000000011010101000000000011110111;
    mem[91] = 162'b000000000011111010000000000000001110000000000011000110000000000011010000111111111111111111111111111101000000111111111100101001000000000100011000000000000001111000;
    mem[92] = 162'b111111111100010001000000000101111011111111111011010111111111111110101110000000000010011011111111111100100000111111111110011001111111111100001011111111111000100010;
    mem[93] = 162'b000000000001000000111111111111000111000000000110010110111111111111011100111111111111111011111111111110100101111111111011011111111111111111001011111111111111111001;
    mem[94] = 162'b000000000001111111000000000000000101111111111011110010000000000010001000000000000000000101000000000010110100111111111001011110000000000110001100000000000100001100;
    mem[95] = 162'b000000000011010101000000000000000110000000000101111010000000000000101111000000000100010100000000000011110011000000000001011010111111111001010110000000000010001100;
    mem[96] = 162'b111111111111110011000000000000000111000000000000001110000000000000000100111111111111110000111111111111100110111111111111101010000000000000001100111111111111110100;
    mem[97] = 162'b000000000000011110111111111111101011111111111111110001111111111111111000111111111111011110111111111111111001111111111111100111111111111111111110111111111111111001;
    mem[98] = 162'b000000000000001111000000000000011001000000000000000011000000000000010110000000000000000001000000000000100100111111111111111111000000000000001111000000000000100001;
    mem[99] = 162'b111111111111101001000000000000000100000000000000001010111111111111111110000000000000010000111111111111111100000000000000001101000000000000000011111111111111110110;
    mem[100] = 162'b000000000000000101000000000000000011111111111111110101000000000000010000000000000000000100000000000000000111000000000000000101111111111111111111000000000000000110;
    mem[101] = 162'b111111111111111101111111111111111001111111111111110010000000000000000111111111111111110111111111111111110111111111111111101000000000000000001100000000000000100100;
    mem[102] = 162'b000000000000001011000000000000000010000000000000001011111111111111101101111111111111110111111111111111110000000000000000001111111111111111111001000000000000000010;
    mem[103] = 162'b111111111111110100000000000000000001111111111111110111000000000000000011111111111111111011111111111111111010111111111111010111111111111111111101000000000000010000;
    mem[104] = 162'b000000000000000001000000000000000000000000000000010010111111111111111011000000000000001010000000000000001100000000000000001100000000000000000100000000000000010101;
    mem[105] = 162'b000000000000000101000000000000001001000000000000000111000000000000001100000000000000001100111111111111111001000000000000000111111111111111100011111111111111111011;
    mem[106] = 162'b000000000000000010000000000000001001000000000000000010111111111111101001111111111111111111111111111111111001111111111111110101111111111111110011111111111111110011;
    mem[107] = 162'b111111111111110111111111111111110101111111111111111100000000000000000001111111111111110010000000000000000000111111111111110111111111111111111000000000000000000000;
    mem[108] = 162'b000000000000010011000000000000001011000000000000000001000000000000001011000000000000000010111111111111111011000000000000001111000000000000000010111111111111111111;
    mem[109] = 162'b111111111111111000111111111111111011000000000000000101000000000000000111000000000000000111000000000000000000111111111111111111111111111111111000111111111111110011;
    mem[110] = 162'b111111111111111011111111111111110110000000000000010010111111111111110011000000000000001101111111111111101100000000000000000000000000000000000001111111111111111100;
    mem[111] = 162'b111111111111110101111111111111111101111111111111110101111111111111110101000000000000000110111111111111101101111111111111101010111111111111111011111111111111111001;
    mem[112] = 162'b000000000000000010000000000000001110111111111111111111000000000000011001000000000000000100000000000000000101111111111111011101111111111111111001000000000000000100;
    mem[113] = 162'b000000000000000110111111111111111010000000000000010110000000000000010001000000000000001010000000000000000110111111111111110101000000000000011000111111111111110111;
    mem[114] = 162'b000000000000001100111111111111111010000000000000000100000000000000000100111111111111111111111111111111111101000000000000000011111111111111111100111111111111110001;
    mem[115] = 162'b111111111111111011000000000000001110000000000000000011111111111111111001000000000000000001111111111111110010000000000000000010111111111111111001111111111111111010;
    mem[116] = 162'b111111111111111111000000000000001111000000000000000000111111111111110101000000000000001001000000000000001011000000000000001101111111111111110110000000000000001000;
    mem[117] = 162'b111111111111111101000000000000001001111111111111101111111111111111110000000000000000000010000000000000001101000000000000000111000000000000001100111111111111101101;
    mem[118] = 162'b000000000000011010000000000000010001000000000000001010000000000000001010000000000000001010000000000000100100000000000000010000000000000000010010111111111111111110;
    mem[119] = 162'b111111111111100001000000000000000111000000000000011000000000000000001010000000000000001010111111111111111111111111111111111110000000000000011001000000000000000111;
    mem[120] = 162'b111111111111111100111111111111110110111111111111111001000000000000000010000000000000001010000000000000001100000000000000001101111111111111110110111111111111110101;
    mem[121] = 162'b111111111111111000000000000000010000111111111111111111000000000000001110111111111111110110000000000000001110000000000000010111000000000000000101000000000000001010;
    mem[122] = 162'b111111111111101010111111111111100011111111111111100010000000000000000011111111111111111110111111111111111111111111111111100110111111111111110110000000000000000101;
    mem[123] = 162'b111111111111111001111111111111110111111111111111110010000000000000000001111111111111111110000000000000000101111111111111111000000000000000000010111111111111111110;
    mem[124] = 162'b111111111111111100111111111111111100000000000000001111111111111111111100111111111111111100111111111111101111000000000000010101000000000000010010000000000000010011;
    mem[125] = 162'b000000000000000001000000000000000011111111111111111111111111111111110100111111111111111111111111111111111100111111111111111111111111111111111010111111111111110011;
    mem[126] = 162'b111111111111111010111111111111100001000000000000001011111111111111111000111111111111111110000000000000000000000000000000010011111111111111111111000000000000000110;
    mem[127] = 162'b111111111111110000000000000000001000111111111111111011000000000000000010000000000000001101111111111111101101000000000000010111000000000000011111000000000000010101;
    mem[128] = 162'b111111111111010111000000000100101001000000000100101110000000000100001010111111111100101111111111111111100000000000000000000111111111111111011001000000000000000111;
    mem[129] = 162'b111111111111111100000000000000000000000000000000001010000000000000001001000000000000011000000000000000000101111111111111111011111111111111101100000000000001111100;
    mem[130] = 162'b000000000000001000000000000000010001000000000000010000111111111111111111111111111111111101111111111111111010111111111111111000111111111111111011111111111111111100;
    mem[131] = 162'b111111111111111001111111111111111100111111111111110100000000000000000100000000000000000001000000000000000101111111111111110001111111111111110101000000000000010000;
    mem[132] = 162'b000000000000000100111111111111110101000000000000000111000000000000000011000000000000010111000000000000000010000000000001000010111111111111110110000000000000001010;
    mem[133] = 162'b111111111111110010111111111111110000000000000000010011000000000000001000000000000000000101000000000000010000111111111111101111111111111111011001000000000001011111;
    mem[134] = 162'b000000000101010111000000000101010100000000000101010100000000000000001000111111111111111111111111111111111101000000000000000111111111111111110100111111111111111001;
    mem[135] = 162'b000000000000011000111111111110110110111111111111111010000000000000000100111111111111100111000000000001101101000000000000011100000000000000001010000000000011011101;
    mem[136] = 162'b111111111111111011111111111111111100111111111111111011111111111111111110111111111111111010000000000000001000000000000000001100000000000000001001000000000000000101;
    mem[137] = 162'b000000000000000101111111111111111011000000000000000100000000000000001001000000000000000011000000000000010011000000000000000101111111111111110101111111111111111001;
    mem[138] = 162'b111111111111111101000000000000000011111111111111110101000000000000000010111111111111110110111111111111111111000000000000000010000000000000000010000000000000000011;
    mem[139] = 162'b000000000000000000111111111111111011111111111111111101111111111111111001000000000000000100000000000000000000000000000000000110111111111111111011000000000000000100;
    mem[140] = 162'b000000000101100010000000000011110111000000000011111100000000000011001000000000000000011001111111111111010010000000000000100010000000000000111100111111111100111011;
    mem[141] = 162'b000000000000000111000000000000000101000000000000000011000000000000000010000000000000000000000000000000000010000000000010101111000000000010000011000000000000111010;
    mem[142] = 162'b000000000010100001000000000011010010000000000101000101000000000000000000111111111111110101111111111111111101000000000000000000000000000000000000111111111111111011;
    mem[143] = 162'b000000000001101000111111111111011101111111111111111000000000000000010100000000000010011110000000000010111111111111111111011101000000000000000101000000000001111010;
    mem[144] = 162'b111111111111110111111111111111111110111111111111111010000000000000000010000000000000000011000000000000000110111111111111111011111111111111111101111111111111111100;
    mem[145] = 162'b111111111111111000111111111111101011111111111111111101000000000000000110000000000000000101111111111111111100111111111111111101000000000000000100111111111111111101;
    mem[146] = 162'b111111111111111000111111111111111110000000000000000010000000000000000110111111111111111111111111111111111101000000000000000001111111111111111000111111111111110010;
    mem[147] = 162'b000000000000000111000000000000000000000000000000000011000000000000000000111111111111111110000000000000000011111111111111111000111111111111111011000000000000000011;
    mem[148] = 162'b000000000000000111000000000000000100000000000000000111000000000000001001111111111111111010000000000000010101000000000000001001000000000000010010000000000000001111;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110100111111111111111100111111111111111000;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule