`include "num_data.v"

module w_rom_14 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000101000110111111110110011010111111111011100000000000000000100010111111111100101100111111111110001111111111111101110110000000000111101111000000000110100011;
    mem[1] = 162'b111111111110100011111111111110110000111111111001111110000000010000010111111111111010101111000000000000100001000000000111111010111111111111101001000000000000011101;
    mem[2] = 162'b111111111101000001111111111111111010000000000010001111111111111111101001000000000010110101000000000011001010111111111101111000111111111110100011111111110111110001;
    mem[3] = 162'b000000000101101010111111111010011101000000001000100110000000010010001101111111110001000101000000001100101110111111111001011101000000010000011111111111111110111110;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b000000000010001011000000001010010000111111110101101110111111110111110111111111111100000100111111111000111000111111111100111111111111111101100010111111111001010100;
    mem[33] = 162'b111111111100011010111111111110011010000000000011101101111111111001111100111111111110111000111111111111001010000000000000010000111111111011111111111111111011000100;
    mem[34] = 162'b000000000000010111111111111111000011111111110110110100000000000000001111111111111110101000000000000011101100000000000001100001000000000000001111111111111101001110;
    mem[35] = 162'b111111111110000101111111111100101111000000000010111110000000001010111110111111111100111000000000000000101100000000000010110001000000000010001011000000000011001010;
    mem[36] = 162'b000000000000000010000000000001001000000000001010101001111111111111110101000000000011010001000000000101000100000000001001010111000000000100010011111111111100010110;
    mem[37] = 162'b111111111110101110111111110110011110000000000010110110111111111100111001111111111111011101111111111101001111000000000001111000000000000010001100000000000110011010;
    mem[38] = 162'b000000000110010001000000001010010110000000000100101101000000000001110101000000000100001111000000000101010001000000000101001000000000000101001010000000000001100001;
    mem[39] = 162'b000000000010110011111111111111101110111111111110010010111111111101000000000000000000111010000000000111100100000000000001010111000000000001110110000000000001000101;
    mem[40] = 162'b000000000010101101000000001011000100000000001001000111000000000000111001000000001100010000000000000111000000000000000001101111000000000101000010000000001000100101;
    mem[41] = 162'b000000000010110000111111111101110110000000000101110010111111111110010110000000000001000010000000000101101001000000000110000100000000001110000001000000000011100100;
    mem[42] = 162'b111111110111011111000000000010111011000000000011010011111111111100110100000000000100100000000000000111010000111111111001101100000000001000001010111111111100111010;
    mem[43] = 162'b000000000100100001000000000110010001000000000010000010111111111001111010000000000011001111111111111110110100000000000111011101000000000000001110111111111111111001;
    mem[44] = 162'b111111110111000111000000000000010100000000000000101000000000000011101000111111111110101101000000000011000000111111111110101101000000000001010000111111111111110000;
    mem[45] = 162'b000000000010011010000000000101010101000000000110111111111111110111010100111111111110100001111111111111000000111111111110101100000000000100000000111111111110101010;
    mem[46] = 162'b111111111101101100111111111101111100000000000101000010111111111111001011111111111100110111000000001001101010111111111100000011000000000001010111111111111100111101;
    mem[47] = 162'b111111111001101100000000001000111110000000000000110111000000000000100011000000000000100110111111111001010100111111111110100001111111111010111100000000000010001110;
    mem[48] = 162'b000000000101010001000000001001100010111111111010110001000000000000100001000000000010101001000000000010110100000000000000010000111111111100110110111111110111000111;
    mem[49] = 162'b000000000001010110111111101101010000000000000011001001111111110110110110111111111010110100111111111010000110111111110111010011111111111010011001000000001000100010;
    mem[50] = 162'b111111111100111100000000000100000001000000000011101001000000000010000000111111111011101011000000000001100010111111111101110101000000000001010001000000001010010011;
    mem[51] = 162'b000000001001111011000000001100110111000000010000011110000000000111001011000000001110111010000000001110111000000000001100010111000000001000100111000000001001000100;
    mem[52] = 162'b000000000111010011000000000101110011000000000110111101000000000110000100000000001101011101000000001001100001000000000011011000000000000000111011000000000110111110;
    mem[53] = 162'b000000000000110110111111111001110111111111111110001000111111111110110001000000000101101110000000000010000111000000000001100101111111111110001100111111111101000011;
    mem[54] = 162'b000000000110010110000000000100110011111111111000110000111111111111001111111111111011000000000000000011111010000000000011011111000000000001111001111111111100010000;
    mem[55] = 162'b111111111111000010111111111111111101000000000001010101111111111101110000111111111011111110111111111011011010111111111111000001000000000001011101000000000110100111;
    mem[56] = 162'b000000000001000100111111111110110011111111111100010101000000000000100100000000000010100111111111111100101100000000000011100010000000000000111010000000000001110011;
    mem[57] = 162'b111111111110110110000000001011011000111111111111011010000000000001111000111111111111100000111111111110001111111111111111011100111111111111111010000000000101001010;
    mem[58] = 162'b000000000011101111000000000101110101111111111100111100111111111011100100111111111111010011000000000011001010000000000101010011000000001001001010111111111101100011;
    mem[59] = 162'b000000000010100101000000001001010010000000000010101111111111111101000111111111111111110110111111111101100001111111111011101000111111111100001111000000001001011111;
    mem[60] = 162'b111111111010100001111111111100001111111111111101011010000000000010111011000000001000001000111111111100011011111111111110000011111111110101101001000000000000001100;
    mem[61] = 162'b000000000010100111000000000001000110000000000101001001000000000000101000000000000010101111111111111110011010111111111101110100000000000100110101111111111110010001;
    mem[62] = 162'b000000001100110000111111111010100000000000000110111100000000000111100011000000000011010110000000000010000011111111111011110001111111111101100100111111111001011110;
    mem[63] = 162'b111111111101110000000000000000000111000000000010010100111111111110111101000000000000010011000000000100000000000000000011101000000000001010101011000000001001110010;
    mem[64] = 162'b111111111100110000111111110110011100000000000010001110000000000110001001111111111101101101111111111110001001000000000100010000111111111110001111000000000100011001;
    mem[65] = 162'b000000000110100000111111111110111001111111111110001010000000000011011101000000000010001110000000000000000011111111111111010111000000000010101010111111111111000000;
    mem[66] = 162'b000000000001001000111111111110111111111111111111111000111111111100001000000000000011110001111111111011000110111111111100011100111111111111101001000000000010111101;
    mem[67] = 162'b111111111100111000111111111111001000111111111000001111111111111110110011000000000010001000000000000000101011000000000001110001111111111110100111000000000110011111;
    mem[68] = 162'b000000000101101001111111111000110010000000000001010011000000000011101111111111111001001101111111111101000000111111111010000010000000000001110000111111111100001010;
    mem[69] = 162'b111111111100010111111111111011011001111111111100111110111111111000001000000000000101010110111111111111001110111111111101011101111111111110100011000000000011111011;
    mem[70] = 162'b000000000000101011000000000011110111000000000001001100111111111101011110000000000110010111111111111011111010000000000001010001000000000000100000111111111111001100;
    mem[71] = 162'b000000000010101011111111111100011011111111111000011101000000000000111010111111111100010011111111111010000011000000000100010100000000000101000111000000000010000011;
    mem[72] = 162'b111111111101001111000000000011010111111111111001100001111111110110010011000000000010110100111111111010101100111111111010111110111111111011100111111111110111001110;
    mem[73] = 162'b111111111101010110111111111100110101111111111110101001000000000000001000000000000011000100111111111110001001000000000001011000000000000000111100111111110111110101;
    mem[74] = 162'b111111111110001011000000000011100001111111111100010010111111111011110010000000000011010110000000000000001100111111111011111011111111111100100111111111111100001111;
    mem[75] = 162'b000000000011001000000000000010100111000000000111011100111111111111111010111111111001100000111111111101011111111111111110001001111111111101100011000000000100011110;
    mem[76] = 162'b000000000111001110000000000101001001000000000100010000000000000111111011111111111100000000000000000011101100000000001001000111000000000100110101000000000001011100;
    mem[77] = 162'b000000000010000000000000000010101100000000000000001001000000000111101100111111111110001110000000000000011011111111111111000110111111110110100011111111110111110011;
    mem[78] = 162'b000000000110000101000000001000001011000000000001100010000000001001100111000000000100101001000000000011010010000000001000010000000000000000000100000000000100110110;
    mem[79] = 162'b000000000000011101000000000001011011111111111110110101000000000000010010111111111101011101000000000001100111111111111111100111000000000011100100000000000101000111;
    mem[80] = 162'b111111111110001100000000000011000001000000000001101100000000000010100001111111111111000011111111111011010100111111111001111010111111111110000011111111111110011011;
    mem[81] = 162'b000000000001000000111111111011111110111111111100100111000000000001010010111111111110011000111111111111011101111111111000111001000000000011001110111111111110010011;
    mem[82] = 162'b000000000011111001000000000001101000000000000001011010000000000010010010000000000000001010000000000001111001111111111100011110000000000101000001000000000000100100;
    mem[83] = 162'b000000000001100011000000000011011011000000000011111111000000000011001100000000000101010110111111111011000011111111111111010110000000000110100110111111111110110100;
    mem[84] = 162'b111111111001001000111111111011110001000000000000010000111111110101001110111111111111110100000000000110000011111111111110011110000000000001011110111111111111100011;
    mem[85] = 162'b000000000011001000000000000011010100111111111010100010000000000110000011111111111100111100111111111110011000000000000000110000000000000010011111111111111111100100;
    mem[86] = 162'b000000000100110111000000000000111101000000000001110010000000000100101001000000000100101001000000000000100011000000001010100011000000000110000011000000000100000000;
    mem[87] = 162'b111111111110011011000000000000100011111111111100000111111111111001000011000000000001001011000000000011001011000000000001101101000000000000000110000000000001011001;
    mem[88] = 162'b111111111111001010000000000001000111000000000010100111000000000001010000111111111011111011000000000000111101111111111011111101111111111111111111000000000100001101;
    mem[89] = 162'b111111111011100010111111111111001001111111111110101110000000000000010001111111111001001110000000000010010001111111111100100101000000000100010111000000000001110001;
    mem[90] = 162'b000000000011001110000000000000100010000000000001111010000000000010011011111111111100100000111111111110100011000000000001011000000000000011111001111111111111001011;
    mem[91] = 162'b111111111111000110000000000100000010111111111110110011000000000010111110111111111111001100000000000010110110000000000100100010000000000011011000000000000110010111;
    mem[92] = 162'b000000000010011100111111111110010000000000000000010001111111111110010010111111111100101000111111111110100011111111111010100110000000000100011001111111111100011001;
    mem[93] = 162'b111111110101001010111111111111101001000000000001111010111111111100011000111111111000001010000000000000110011000000000000000000000000000010011111000000000010010100;
    mem[94] = 162'b111111111010001010000000000001001100000000000001010100111111110111010111111111111001100011000000000010111010111111111100011011000000000001101111000000000001011001;
    mem[95] = 162'b111111111110110111111111111100110011111111111101111110111111111101001000000000000010000010000000000100001100000000000101000011111111111111110010000000000010101011;
    mem[96] = 162'b000000000000010100111111111111111000000000000000010001000000000000010001111111111111111111000000000000011000111111111111110011111111111111111001000000000000000001;
    mem[97] = 162'b000000000000001000111111111111111001000000000000001010000000000000001011000000000000011001111111111111110001000000000000010111111111111111101011000000000000010001;
    mem[98] = 162'b000000000000001100111111111111111111111111111111110001111111111111111110000000000000010000111111111111111111000000000000000101000000000000000111000000000000000011;
    mem[99] = 162'b000000000000001010000000000000000101000000000000011001111111111111111000111111111111111011000000000000000100111111111111101111000000000000000000000000000000000011;
    mem[100] = 162'b000000000000001101000000000000001111000000000000000101111111111111111000111111111111110101000000000000000000000000000000000010111111111111111001111111111111111100;
    mem[101] = 162'b000000000000101011000000000000010111000000000000011110000000000000000010000000000000000001000000000000000010000000000000010101000000000000000101111111111111111111;
    mem[102] = 162'b000000000000000111000000000000001101111111111111111001111111111111110001111111111111111011000000000000000001000000000000000000000000000000000110000000000000000010;
    mem[103] = 162'b111111111111101110000000000000000101111111111111111001000000000000000011000000000000001110111111111111111111111111111111101111000000000000000010000000000000001000;
    mem[104] = 162'b111111111111111010000000000000001101000000000000001100000000000000001110000000000000001000000000000000001111000000000000001000000000000000001011000000000000000011;
    mem[105] = 162'b111111111111110010111111111111110110000000000000010001000000000000011000111111111111111000111111111111111010111111111111111111000000000000000111111111111111110010;
    mem[106] = 162'b000000000000000111000000000000001001000000000000001100000000000000000100000000000000010001000000000000001100000000000000000110111111111111111000000000000000011110;
    mem[107] = 162'b111111111111111000111111111111110010111111111111111010111111111111101010111111111111111010111111111111100110111111111111110110000000000000010110111111111111111110;
    mem[108] = 162'b000000000000000001000000000000011100000000000000000011000000000000010010000000000000001010000000000000010101000000000000001011000000000000010000111111111111111100;
    mem[109] = 162'b000000000000010110000000000000001001000000000000000011000000000000001010000000000000001001000000000000000001111111111111110111000000000000000110000000000000001111;
    mem[110] = 162'b000000000000000110000000000000001111000000000000000100111111111111110100000000000000000010111111111111101010000000000000001101111111111111110001000000000000010101;
    mem[111] = 162'b000000000000001000000000000000000110000000000000001001111111111111111010000000000000010010111111111111110000111111111111111000000000000000000110000000000000001110;
    mem[112] = 162'b000000000000011110000000000000011001000000000000101000000000000000100111000000000000000011000000000000011001000000000000010100111111111111111111000000000000011001;
    mem[113] = 162'b000000000000010011000000000000000000000000000000000111000000000000000101000000000000010011111111111111011010000000000000100011111111111111111101000000000000001011;
    mem[114] = 162'b000000000000000011111111111111111011000000000000000100111111111111111100111111111111111011000000000000000110000000000000000111111111111111110011111111111111111100;
    mem[115] = 162'b111111111111110010111111111111111101000000000000000110111111111111101001000000000000000010000000000000001000000000000000011001000000000000010110000000000000000111;
    mem[116] = 162'b111111111111101101111111111111111100000000000000000000111111111111111011111111111111100100000000000000000111111111111111110010111111111111111100111111111111110010;
    mem[117] = 162'b111111111111110101000000000000000100111111111111101110000000000000010001111111111111111010111111111111111100000000000000000111000000000000000100000000000000000101;
    mem[118] = 162'b000000000000101100000000000000000011000000000000001011000000000000001110111111111111101111111111111111111001000000000000000101000000000000001000000000000000001111;
    mem[119] = 162'b000000000000001001000000000000000010111111111111111001111111111111111110111111111111111011000000000000011011111111111111111110111111111111111010000000000000000011;
    mem[120] = 162'b000000000000001100111111111111110110000000000000000101000000000000001110000000000000001011000000000000000110000000000000001100000000000000001000111111111111101111;
    mem[121] = 162'b000000000000011001000000000000001001000000000000110111111111111111110001000000000000000111000000000000011100111111111111110011000000000000101011000000000000101110;
    mem[122] = 162'b111111111111110100000000000000010011111111111111111000000000000000000100000000000000001010000000000000000010111111111111111110000000000000000010000000000000010010;
    mem[123] = 162'b000000000000000000111111111111110011000000000000001100111111111111110110000000000000001101111111111111111100111111111111110001111111111111110000111111111111101011;
    mem[124] = 162'b111111111111110001000000000000000100000000000000001100000000000000001110111111111111111101000000000000001011111111111111111010000000000000001011000000000000010100;
    mem[125] = 162'b111111111111100111111111111111110110111111111111101100111111111111100010111111111111101010111111111111110111111111111111111101000000000000010001000000000000001101;
    mem[126] = 162'b000000000000010101111111111111111011111111111111111101111111111111111010000000000000000000111111111111110101000000000000000101111111111111110110000000000000000111;
    mem[127] = 162'b111111111111111000111111111111111001111111111111111100111111111111111000111111111111101011111111111111111001111111111111110001111111111111110010111111111111110000;
    mem[128] = 162'b000000000000100000000000000100111011000000000101010101000000000100010010000000000000000001111111111111111011000000000000100001000000000000001001000000000000100100;
    mem[129] = 162'b000000000000000000000000000000000011000000000000001010000000000000000111000000000000000110111111111111111110000000000000101000000000000000001101111111111110111110;
    mem[130] = 162'b000000000000000110000000000000000010000000000000000110000000000000000101000000000000000101000000000000000010000000000000000000111111111111110001111111111111111011;
    mem[131] = 162'b000000000000000010111111111111111110111111111111111010000000000000000000000000000000000100000000000000000110000000000000000101000000000000001100000000000000010100;
    mem[132] = 162'b000000000000101111000000000000001100000000000000000001000000000000001111111111111111010000000000000000000000000000000000011011111111111111010011000000000000001011;
    mem[133] = 162'b000000000000000010000000000000000000000000000000010010000000000000001000000000000000000110111111111111111001000000000000010010111111111111101010111111111111100011;
    mem[134] = 162'b000000000101011011000000000101001110000000000001111000000000000000001101000000000000000001111111111111111111111111111111111100111111111111110001111111111111111011;
    mem[135] = 162'b000000000000010101000000000010000001000000000000111100111111111111101100000000000000101000000000000010000101111111111111011001111111111111100111000000000001110111;
    mem[136] = 162'b111111111111101111111111111111101111111111111111110000111111111111111000111111111111110101000000000000010101000000000000000001000000000000000000111111111111111100;
    mem[137] = 162'b000000000000001101000000000000001001000000000000001001111111111111111000111111111111111111000000000000000101111111111111111001111111111111110110111111111111111100;
    mem[138] = 162'b000000000000000101111111111111111100111111111111111101111111111111111111111111111111111011000000000000001100111111111111111100111111111111111110000000000000001100;
    mem[139] = 162'b111111111111111111000000000000001111111111111111111111111111111111111111000000000000001001000000000000000100111111111111111011111111111111111110000000000000001110;
    mem[140] = 162'b000000000001011011000000000001101101000000000101010001000000000011101101000000000000011010111111111111111100111111111111101111000000000000000011111111111101011100;
    mem[141] = 162'b111111111111111111000000000000000000111111111111111110111111111111111101111111111111111110000000000000000111000000000011000000000000000001011111000000000000110000;
    mem[142] = 162'b000000000011110100000000000100000110000000000100110000000000000000000001111111111111110111111111111111110010111111111111111111000000000000000001111111111111111101;
    mem[143] = 162'b000000000011010000111111111111100000000000000000000110111111111111011101000000000001011100111111111111001001000000000001011111111111111111011100000000000001100100;
    mem[144] = 162'b111111111111111010111111111111111101111111111111111110111111111111110111111111111111110010111111111111111000111111111111110111111111111111110010111111111111111011;
    mem[145] = 162'b000000000000000110111111111111111000111111111111110111111111111111111010111111111111110011111111111111110110111111111111111101000000000000001101000000000000000010;
    mem[146] = 162'b000000000000000100111111111111111111111111111111111011111111111111111011000000000000000010000000000000001001111111111111111001111111111111100111111111111111110111;
    mem[147] = 162'b111111111111111011000000000000000000000000000000000001000000000000000000000000000000000011000000000000000111111111111111111111111111111111110110000000000000000011;
    mem[148] = 162'b111111111111111110000000000000000110000000000000001111000000000000001000111111111111111001000000000000001100000000000000000110000000000000000000000000000000001000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110111000000000000000100111111111111111110;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule