`include "num_data.v"

module w_rom_27 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000011101011000000000100110001000000000010100001000000000011001111000000000011010010000000001000001001111111111110101000111111111101010001111111111110000111;
    mem[1] = 162'b000000011000001001111111111010110010000000000110100111111111111100101100000000010100101011111111110110000010111111111111011001000000000001001000000000000111110100;
    mem[2] = 162'b111111111111101101111111111111111110111111111101110101111111111111001001111111111100100111111111111101111010111111111110100111111111111101111111111111111110111100;
    mem[3] = 162'b111111110001110001000000000000110100111111110001110100000000010111000011000000000011011010111111111111011100111111110100011010111111111110100100000000000001111000;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111111001001111111111100010111111111111111101001111111111110110001000000000010100011111111111111011101000000000100011010111111111111010111111111111101001110;
    mem[33] = 162'b111111110110111100000000000100011011000000000101111110111111111111000011000000000010011011000000000000000100111111111010011010000000000100011100111111111100101101;
    mem[34] = 162'b111111111010010000111111111100111111111111111101001111111111111100110100000000000001011011000000000011100000111111111001111000000000000001101000111111111001110000;
    mem[35] = 162'b000000000000001110000000000001110010000000001000000100000000000100110111111111111010000001000000000001001110111111110101001011111111110110101110111111111011111101;
    mem[36] = 162'b000000000001001001000000000101001111000000001000100010000000000010011100000000000011110100000000000101110101000000000000001110111111111100110011111111111001001100;
    mem[37] = 162'b111111111100101101000000000101110011000000000010111001000000000001101010111111111110011010000000000001001011111111110110000110111111111110011101111111111111000011;
    mem[38] = 162'b000000001001010011000000000000100100000000001001100001000000000100011011000000000110110101000000000111111000000000000101000111111111111110001000111111111101011101;
    mem[39] = 162'b000000000010001100000000000101111010000000000100000101111111111110001100000000000100000011000000000000110001111111111110101100000000000001111111111111111011111111;
    mem[40] = 162'b000000000101110001000000001001000111000000001010000111000000000101001101000000000001111011000000000100111010111111111011011000111111111101001000111111111111100001;
    mem[41] = 162'b000000000101011101000000000011011011000000000000111000111111111001010000111111111111100101111111111110001110111111111100001011111111111011001010000000000011010000;
    mem[42] = 162'b111111111010100010111111111110000000000000000110000010000000000110000001000000000110000111111111110110010101111111111001010000000000000001000001111111110110101111;
    mem[43] = 162'b000000000111110101000000000101111101000000000111100011000000000100011011000000000011000110000000000100001001111111110111010100111111110000100001000000000001011101;
    mem[44] = 162'b000000000010101000111111111101011111000000000001001100111111111111111101000000000000010110000000000100001101111111111010101011000000000000011110000000000000010000;
    mem[45] = 162'b111111111110001100000000000100011000111111111111100001111111111101001101111111111000101101000000000001111001111111111011000111000000000000111011111111110111000101;
    mem[46] = 162'b111111111101000000000000000010101100000000001001101000111111111011011001000000000000100101000000000000000010111111111111010010000000000100001111111111111100101010;
    mem[47] = 162'b111111111111010001111111111011101111111111111011000000000000000011010010000000000001101011000000001011000000111111111101000010000000000000110101111111111111110000;
    mem[48] = 162'b111111110111101000000000000010000001000000000101010011111111111110100000111111111110111000000000000000110001111111110110010111000000000110101101111111110001001101;
    mem[49] = 162'b111111111111111011111111110110111111111111110000010111000000000001010011111111111101010110111111111111110101000000000101010001111111111010111110000000000101001010;
    mem[50] = 162'b111111111111111101000000000110000000111111111110101010111111111011100111111111111110110111000000000000001101000000000001000011000000000001111100000000000000001011;
    mem[51] = 162'b000000001011111011000000001111011011000000001110010010000000001000101010000000000101111001000000001000100011000000000110101010111111111111101001000000000011101110;
    mem[52] = 162'b000000000110010100000000001011100100000000000111110011000000000011010001000000000101101000000000001000011110111111111011101011111111111100101011111111110011000010;
    mem[53] = 162'b000000000001000101000000001011111000111111111100110010000000000011100100000000001010000111000000000001101001111111111100100110111111111001010101000000000000010010;
    mem[54] = 162'b000000001000110010000000000100001111111111111010010100111111111110110000111111111111010110111111111100011011000000000011011000111111111111000101111111111101110010;
    mem[55] = 162'b111111111100101101000000000001000110111111111101100101000000000001010000111111111111110101111111111111011010111111111100001010111111111111101011111111111011010101;
    mem[56] = 162'b111111111110000010111111111010110011000000000101000100111111111100100000111111111111001110111111111111100000111111111111101001000000000100110010111111111101001110;
    mem[57] = 162'b111111110101010010000000000110010111111111111001111100000000000000010001111111111111100101000000000000110001000000000010011101111111111010001101000000001001100110;
    mem[58] = 162'b000000001001010011000000000001010000000000000100000100111111111111110100000000000101001111000000001000000110000000000101010100111111110110000110111111110010011101;
    mem[59] = 162'b111111111101011111000000000100100010111111111101001011111111110001101000111111111110100000111111111110010011000000000001110001111111110101000111111111111110001111;
    mem[60] = 162'b000000000101100010111111111101011001000000000000011101000000000010100010000000000001111101111111111111111111111111111101110111000000000000100111000000000001111000;
    mem[61] = 162'b000000000010010110000000000110101001111111111000111100000000000100010000111111111011100010111111111011110000000000000010100001111111111111101000111111111110010110;
    mem[62] = 162'b000000000001111011000000000011100010000000001100010010111111111110011111111111111111001000111111111011111101000000000000101110111111110111000100000000000010011011;
    mem[63] = 162'b000000001010101001000000000101111101000000000001100111000000000010101010000000000001110001000000000101011001111111111110000001111111111101011111000000000000001100;
    mem[64] = 162'b111111110110111001111111110101001001111111111010011110111111111011111110000000000011001110111111111110010110000000000100000001111111111111101110111111111001110101;
    mem[65] = 162'b000000000000101001000000000001110010000000000000000010000000000010011001000000000001000110000000000001000010111111111111100000000000000101011011000000000110111100;
    mem[66] = 162'b000000000010110000111111111010000001111111111110001011111111111110010010000000000000001010111111111011010001000000000100011111000000000000100011000000000000110100;
    mem[67] = 162'b111111111111110010111111111111010010111111111010000111111111111110010100000000000000101100000000000000011110000000000011010101111111111111011100111111110111001101;
    mem[68] = 162'b000000000001001011111111111110111001111111111110110011000000000000000100000000000001011110111111111110011111111111111111110001000000000000001100000000000000000100;
    mem[69] = 162'b000000000101100010111111111101111110000000000010111110000000000000100000111111111001111001111111111110010001111111111110110000000000000011100111000000000110001110;
    mem[70] = 162'b111111111100111011000000000011101011000000000011011100000000000010000111000000000000111100000000000001110100111111111110100100000000000100010101000000001011010101;
    mem[71] = 162'b000000000100110101000000000001101111000000000000010011000000000100011110111111111011010000000000000100111110111111111111011011000000000011000001000000000100001100;
    mem[72] = 162'b000000000100110000000000000011100100111111111111001110111111111111000011111111111101111011000000000100010110111111111101101110111111111100110000111111111101110010;
    mem[73] = 162'b111111111110001010000000000000011101111111111111010110111111111011100010111111111111100001000000000001110111000000001001100111111111111110001011000000000000000000;
    mem[74] = 162'b000000000000111100111111111001111011000000000010000011000000000011000010000000000010010000000000000011100111111111111111010111111111110011110110111111111011010101;
    mem[75] = 162'b000000000000001111000000000110110000000000000100111110111111111110000001000000000100001110111111111100101100000000000001000010000000000100011101111111111100110110;
    mem[76] = 162'b000000000001100101000000000011000110000000000001011001111111111110110001000000000011011001000000000101000010000000000011110011000000000100010000000000001000001001;
    mem[77] = 162'b000000000000101010111111111111111010111111111101011010000000000010101110000000000001111011000000000011011111111111111100110110000000000011110000000000000000010111;
    mem[78] = 162'b000000000010101101000000000011111011111111111111100010000000000001000111111111111111100010000000000110100110000000001000001011000000000010101011000000000011011101;
    mem[79] = 162'b111111111010001111000000000001110101000000000100111111000000000010011110111111111111000001000000000100011010000000000001111100111111111010101111111111111101001011;
    mem[80] = 162'b000000000011001000111111111110111110111111111111010100000000000010101011000000000000110101000000000000100100111111111110010110111111111010011110111111111100011100;
    mem[81] = 162'b111111111000011101000000000000100010000000000010011110000000000000100110111111111100111101000000000100000101000000000000011101111111111110101001111111111100001010;
    mem[82] = 162'b000000000010101101000000000101100001111111111011001110111111111101111010000000000101111111111111111100111100000000000110010101000000000010010100000000000000100110;
    mem[83] = 162'b000000000001010010111111111110101100000000000100111010111111111101001010111111111011101111000000000000010011000000001001000100000000000101111111000000000001010011;
    mem[84] = 162'b111111111111000011111111111110010000000000000011101000000000000100001001111111111110011001000000000100010100000000000100001010000000000011001001111111111110011001;
    mem[85] = 162'b000000000000000100111111111111011100111111111010010001111111111001110010000000001001010011000000000011000010000000000000101001111111111010101111000000000011100000;
    mem[86] = 162'b111111111111111011000000000010000001000000000001001110000000000011010101000000000001001101000000000011001011000000000111011111000000000110011011000000000111011000;
    mem[87] = 162'b111111111010001001000000000010011000000000000011110000111111111100101111111111111000100101000000000000000010111111111110001111000000000010001110111111111011001010;
    mem[88] = 162'b000000000011010110111111111111110011000000000001000101000000000100010101111111111011111101111111111001001011111111111111100001111111111110111100111111111100000111;
    mem[89] = 162'b111111111011110000000000000001011000000000000000100100111111111111010011000000000011100001000000000000000110111111111101001101000000000000101110111111111011100001;
    mem[90] = 162'b111111111111111011000000000000111000000000000111100110111111111011100001111111111101100010000000000000010000111111110110000110111111111011101100000000000111110001;
    mem[91] = 162'b111111111111001101000000000010110010111111111100000000000000000000110101000000000001100110000000000001000011000000000100001110000000001001111011000000001001011011;
    mem[92] = 162'b111111111000011100000000000001010010000000000001010011000000000111110011111111111011000011111111111111110000111111111101010111000000000010100100000000000000110100;
    mem[93] = 162'b111111111101010110000000000000100001000000000010000001000000000010011001111111111100110110000000000000001111000000000001001010000000000011111110111111111111111110;
    mem[94] = 162'b000000000011100100111111111100000110111111111110000011111111111011000011111111111110101111111111111110111000000000000010111001111111111011100110000000000010001010;
    mem[95] = 162'b111111111101101111111111111000101001111111111101000101111111111111111111000000000011100001000000000110111110111111111100111011111111111110101001000000000011101011;
    mem[96] = 162'b111111111101111000111111111110110101111111111111101000111111111111010001000000000000011100000000000010010110111111111110110100111111111100001001111111111101111100;
    mem[97] = 162'b000000000100000000000000000000100111111111111101110010111111111101011100000000000000010110111111111111000001111111111110111100000000000000101101111111111100001010;
    mem[98] = 162'b000000000000011100000000000000001101111111111111111001111111111111011011111111111110111101111111111110000101000000000010001001000000000000001100000000000000110000;
    mem[99] = 162'b000000000010011010111111111101100000000000000010000111111111111110000101111111111001001111111111111100111111111111111001011100111111110110100011000000000001001000;
    mem[100] = 162'b000000000110001011000000000110011001000000001000111000000000000100010010000000000101011110000000000001010011000000000100111011111111111111111010111111111101000000;
    mem[101] = 162'b000000000000110110000000000001010001111111111100110101111111111110110111000000000000001000000000000001100000000000000010000110111111111111111001000000000000111110;
    mem[102] = 162'b111111111100001010111111111111011110000000000001111110111111111111010110000000000000111010111111111111110010111111111101110100111111111011001110111111111110000000;
    mem[103] = 162'b000000000001000001000000000000010111000000000010000110000000000010110110111111111111100110111111111110100101111111111111011110000000000010100011111111111010110011;
    mem[104] = 162'b000000000000111010111111111101100000111111111111000111111111111101110011111111111111110110111111111010100101000000000001100101000000000001010101000000000010001111;
    mem[105] = 162'b000000000001000000000000000010101001111111111101010000111111111110010100111111111101101101000000000010110110111111111110001110111111111110011111111111111010100000;
    mem[106] = 162'b111111111101110010111111111101110010111111111000000001000000000000010001111111111111111101111111111100010101111111111010010000111111111101100101111111111011110110;
    mem[107] = 162'b111111111110000011000000000010001000000000000000110110111111111111111000000000000000101101111111111110111001111111111111100001111111111011010100111111111110010011;
    mem[108] = 162'b000000000010101010000000000000100111111111111110101010000000000001010011111111111111110010111111111110010001111111111100010001000000000010001001111111111101111011;
    mem[109] = 162'b000000000011000111111111111111100101000000000000010110111111111100100110111111111101010000000000000000001011111111111110110000111111111101100000000000000000111101;
    mem[110] = 162'b111111111001000101111111111111001000000000000010001110111111111110110000000000000001000111000000000000001001000000000000010101000000000000101100111111111100111101;
    mem[111] = 162'b111111111101001011111111111110001110111111111011010011111111111111010110111111111111100111111111111111100101111111111111101100000000000000011001111111111110000111;
    mem[112] = 162'b000000001100101101000000001101100001000000001011110011000000010010011100000000001100001011000000001011101111000000000110100010111111111101111111000000000101000101;
    mem[113] = 162'b000000000000110001111111110111001101111111111110011110000000000001010011000000000000011100000000000001010000111111111110111010111111111111111100111111111101111111;
    mem[114] = 162'b000000000100011011000000000100010000000000000011111100111111111011111001111111111011011011111111111011111100000000000010001001000000000000101111000000000000111010;
    mem[115] = 162'b111111111011101000000000000000100010000000000001000000111111111011111000000000000000111111000000000001100100000000000000011001111111111111100101111111111101111011;
    mem[116] = 162'b111111111110001100111111111100000001000000000001001010000000000001000000000000000000000001111111111100110010000000000001001110111111111111111110111111111100100111;
    mem[117] = 162'b000000000000100010000000000000010000111111111100110100000000000000011101111111111101100000111111111110111110111111111111111100111111111110101101000000000000101011;
    mem[118] = 162'b000000000010011010000000000000100011111111111111010010000000000000011001111111111110000011111111111111100011000000000000101010111111111101100111111111111111000101;
    mem[119] = 162'b000000000001111110000000000001010101111111111111110000000000000000011110111111111110010111000000000001110111000000000010010001000000000011010010000000000011011100;
    mem[120] = 162'b000000000001010110000000000000011101111111111011101001111111111100000101111111111111010100111111111111000111111111111101001100000000000000000000111111111111101001;
    mem[121] = 162'b000000001000011111000000000111111101000000001001011100000000001110100010000000001101110011000000001011101000000000000101001100111111111110100011111111111111010011;
    mem[122] = 162'b000000000001001010111111111111001000111111111110011100000000000001110111000000000000111011111111111101001111111111111110111101111111111110100101111111111110011000;
    mem[123] = 162'b000000000001110101111111111111100011000000000000101111111111111110101111111111111111010000111111111111000011000000000001001110111111111110011010111111110111001000;
    mem[124] = 162'b000000000001111100111111111101100001111111111101101100111111111100111000111111111111101011000000000010111000000000000000011000000000000001011001111111111010101100;
    mem[125] = 162'b000000000010011101111111111001010101111111101010101000000000000000010001111111111001111111111111110101110000111111111111011110000000000001110111111111111101111101;
    mem[126] = 162'b000000000000100100000000000000110011111111111111010101000000000010000001000000000000000011000000000000001100000000000000110011111111111101100010111111111011111000;
    mem[127] = 162'b000000000001110000000000000010001000111111111110100011000000000100010011111111111111111011000000000001010110000000000000000110111111111111001111111111111110011110;
    mem[128] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[129] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[130] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[131] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[132] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[133] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[134] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[135] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[136] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[137] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[138] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[139] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[140] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[141] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[142] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[143] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[144] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[145] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[146] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[147] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[148] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule