`include "num_data.v"

module w_rom_8 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b111111111001001110111111111111100100111111111000011101000000000111111010111111111010111001111111111001010001000000000001010011111111110110101011000000000101000101;
    mem[1] = 162'b000000000011001011111111111100000010000000001110011000111111111101101111111111110100111010000000000010110010000000000110111101111111110001110101000000000010100010;
    mem[2] = 162'b111111111011010011000000000011000110000000000010110011111111111010110001111111111110000101000000000100000001000000000010000011111111110011000110111111111010010100;
    mem[3] = 162'b000000001000011101111111111000110110111111111111011110111111111000100101000000001001111101000000000101001110111111111100001000111111010110001001111111100110011011;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b000000000011110011000000000010101100111111111100010001000000000001101101000000001000001011111111111010111101111111111110111110111111111001011010000000000100100001;
    mem[33] = 162'b111111111011011100111111110101100101000000000100000000111111111111100100111111111001000000000000001000010110111111111100111000000000000001101010111111111010010011;
    mem[34] = 162'b111111111100000110111111111011111000111111111000000101000000000011111011000000000001101011111111111101110100000000000110101010111111111000110110111111111101101000;
    mem[35] = 162'b111111111110000100111111111111110000111111111101010110000000001000011010000000000110000000000000000100100110000000000111110010000000000000101000111111111101100010;
    mem[36] = 162'b000000000001011010000000000001000101111111111111001110111111111001101101111111111111101110000000001101110110000000000000100011000000000001001110000000000000101100;
    mem[37] = 162'b111111111010111111111111111000111000111111111111100001000000000100101111000000000010110100111111111010111000000000000100001011111111111100010101111111111111110010;
    mem[38] = 162'b000000000110011011111111111001101010000000000011100000000000000110010001000000000101001111000000000111000111000000000001100000111111111111010000000000001000010101;
    mem[39] = 162'b000000001000100010000000000101110010111111111100111100000000000111000010000000000000101101111111111011100111000000000000110011000000000010000010000000000001011001;
    mem[40] = 162'b000000000110001010000000000100100001000000000111011100111111111100001110000000001000011101000000001001001001111111111010001001111111111011110101111111111010101010;
    mem[41] = 162'b111111111110010011111111111001011011000000000011110001111111111001100110000000000001101100000000001001010101000000000011001011000000000010010110000000000110000101;
    mem[42] = 162'b000000000000110011000000000001011001000000000010010110111111111101010100000000000100000100111111111010101010111111110110001111111111111101100101000000000101111100;
    mem[43] = 162'b000000000011111111111111111101001100111111111110010100000000000010111100111111111111011011000000000101110011000000000001111110111111111001100101000000000001101011;
    mem[44] = 162'b111111111011000010000000000111100100000000000000011111000000001001000000111111111111011101111111111100011000000000000001001100111111111110010000111111111101111111;
    mem[45] = 162'b111111111100010010000000000100010111111111111100111110000000000000110100111111111010111111000000001011000011111111111000010011111111111110110111111111110110100010;
    mem[46] = 162'b000000000001001001000000000010111111111111111100110000000000000100011001111111110111011100000000000011111001111111110110100100000000000101110101111111111000100101;
    mem[47] = 162'b111111111010001010000000000111111000111111111011011101111111111011101111000000000000010100111111111001000111111111111010111010000000000111101000111111111010111001;
    mem[48] = 162'b111111111011110100000000000110000100111111110111101010111111111101001011111111111101100001000000000000101110111111111111111000000000000110010000111111110011011111;
    mem[49] = 162'b000000000100001110111111111110110011000000000000101000000000001011101011111111111100101110111111110100000000000000000101001001111111111000111110111111111001011010;
    mem[50] = 162'b111111111110100011111111111010010110000000000100110000000000000001100010111111111011111100000000000101100000111111111110000100111111111100101101000000000001100100;
    mem[51] = 162'b000000000100000011000000000000110101000000000100000100000000001000000000000000000011110011000000001001010001111111111110100011000000000010101000000000000101010111;
    mem[52] = 162'b000000000000101010111111111110101000000000000100101001000000000100100010000000000001010001000000000110111000000000000100000011000000000000101010000000001101011100;
    mem[53] = 162'b111111111111110000111111111101101110111111111011001001111111111101100101111111111110101011111111111111010011000000000010010011111111111110100010111111111110111100;
    mem[54] = 162'b111111111100111101000000000010101110111111110101101111000000000011100110000000000000111000111111111010100010000000000011110000000000000011010111111111111111101100;
    mem[55] = 162'b111111111110100101111111111011101111000000000011101111000000000001011011000000000101101001000000001001001111000000000101100100000000000001111110111111111111111110;
    mem[56] = 162'b111111111111001110000000000110101100111111111100011011000000000110001100111111111111100110111111111000101110000000000010000110111111111100110110000000000001000110;
    mem[57] = 162'b000000000010110001111111111100110010111111111100110101000000000111110100111111111000111011000000000000010111000000000101100110000000000011100111111111111111011100;
    mem[58] = 162'b000000000011011001111111110111001001000000000100111101000000000111001010111111111111101001000000000111010011111111111010110000000000000001111001111111111110110100;
    mem[59] = 162'b000000001000001111111111111110101011111111111011100110000000000101110111000000000110100101111111111010111000000000000111000000111111111011100100111111111110011110;
    mem[60] = 162'b000000000000011110111111111111101000111111111010110100000000000001000000000000000010000110111111110101110000111111111111111110000000000010110111111111111000110100;
    mem[61] = 162'b000000000010100001111111111011000100000000000001000010000000000011100111111111111000111001000000000000000101111111111010101100000000000010001111111111111100110111;
    mem[62] = 162'b000000000110100101111111111000000111111111111100000001000000000101000011000000000111010010111111111111111100111111111101001011111111111101010000000000000001010000;
    mem[63] = 162'b000000000010000111111111111001110011000000000001111111000000001000101000111111111101011111000000000110011010111111111100111101000000000110000010000000000110010011;
    mem[64] = 162'b111111111100001100000000000000101111111111111011011100111111111111110001000000000001010110000000000010111011111111111111100111000000000010001100111111111111101110;
    mem[65] = 162'b000000000001110011111111111101111001000000000000011010111111111101000110111111111111111100111111111101000101000000000001010100000000000101011111111111111101100100;
    mem[66] = 162'b111111111110010011111111111011101000111111111100101110000000000100110001111111111001001010111111111101001111000000000101001011111111111110011011111111111100010101;
    mem[67] = 162'b000000000000000110111111111110100110000000000000010111000000000010100101000000000010111011111111111011001110111111111111101111111111111111000110000000000000011011;
    mem[68] = 162'b000000000010110011111111111011000111111111111110010110111111110111100101111111111111001000111111111010001001111111111110111010111111111010101111000000000000001111;
    mem[69] = 162'b000000000000011000000000000001000001000000000001110001111111111101100110111111111010101101000000000001010011000000000101101110111111111111000010000000000000111010;
    mem[70] = 162'b111111111101100011000000000011011001000000000011001111111111111101010110000000000000110001111111111100001000111111111011010111111111111101001111111111111111110111;
    mem[71] = 162'b000000000011000001111111111111000100111111111110111101111111111101100000000000000010010111111111111110001010111111111110011110000000000000011111111111111101110011;
    mem[72] = 162'b111111111100111001111111111110100101111111111011001111111111111001100001000000000000100011111111111100111010111111111000100010000000000000111110111111111100011000;
    mem[73] = 162'b111111111110101000111111110101011001111111111000100011111111111111110110111111111111110000111111111000111000000000000100011111111111111101011001111111111111000010;
    mem[74] = 162'b111111111101001010111111111111110010111111111001011000111111111101111000111111111101000111111111111011110100111111111110110010111111111101100110111111111011001010;
    mem[75] = 162'b111111111110010100000000000100111001111111111111110101111111111110100100111111111100000011000000000000011001000000000000101110111111111110111001111111111000100100;
    mem[76] = 162'b000000000110010010000000000101000011000000000100001101000000000101010000000000000011110111000000000101111011000000000010110000000000000011010001000000000101101100;
    mem[77] = 162'b000000000111011000000000000110001011111111111011010001111111111010101000111111111011000110111111111101111001000000000000001100111111111110001100111111110110110000;
    mem[78] = 162'b000000000011010100000000000101100110000000000111001111000000000110101000000000000110011010000000000011001000000000000110011110000000000001101100111111111101001000;
    mem[79] = 162'b111111111111111011000000000011001110000000000011000000111111111111001010000000000010101100000000000000011010000000000000101000000000000100010011000000000101100000;
    mem[80] = 162'b000000000000110111111111111001101110000000000000111110111111111011110000111111111100000100111111111001000000111111111010000001111111111100000011000000000001010111;
    mem[81] = 162'b111111111101000000000000000010101010111111111101110010000000000100001001111111111111001100111111111101000111111111111100000010111111111110101011111111111011000011;
    mem[82] = 162'b111111111111001011000000000011111111000000000100100010000000000010011101000000000000010001111111111101100000111111111011101011000000000010111101111111111111100000;
    mem[83] = 162'b111111111110011111000000000010101000000000000001100000111111111010001111000000000000100101000000000011110111000000000010001111000000000100101111000000000010011010;
    mem[84] = 162'b111111111100010001000000000010011111111111111010011101000000000001000001111111111110101001111111111110011111111111111110010010111111111110101011000000000001111011;
    mem[85] = 162'b111111111110110111000000000000010000111111111111000011000000000100001101000000000110010100111111111100111010111111111111110001000000000101100001000000000010110110;
    mem[86] = 162'b000000001000100100111111111100111101000000000001001101000000000011000110000000000101101111000000001010001011000000001000000101000000001001001010000000000101101000;
    mem[87] = 162'b000000000010001010111111111101011101111111111111001010000000000001101011111111111111100010000000000001001010111111111110010011111111111100110011000000000001000001;
    mem[88] = 162'b111111111010111010111111110110010011111111111011001000000000000000011011111111111010011101000000000001000101111111111011101111111111111110111011000000000000010100;
    mem[89] = 162'b111111111110111100111111111111111111000000000001000001111111111110101001111111111101100011111111111111000001111111111100100101111111111001000011111111110110101011;
    mem[90] = 162'b000000000000111001111111111110010001000000000101001110111111111110101010111111111100011111111111111111111100111111111010110101000000000001101011000000000010011001;
    mem[91] = 162'b111111111110101101111111111100000100111111111111011000000000000001101111000000000010000101000000000011000101000000000001101101000000000011010010000000000010101100;
    mem[92] = 162'b000000000001010101000000000011001111000000000010110110111111111111001010000000000000110001111111111010111010111111111010001011111111111111011010111111111110010011;
    mem[93] = 162'b000000000000111101111111111011101101111111111010101001111111111110011101000000000010111101111111111110100010111111111000111011111111111100011110000000000011010110;
    mem[94] = 162'b111111110111010000000000000100101000111111111101111110111111111111000101000000000010100010000000000001011000000000000010111001111111111100010111000000000010001110;
    mem[95] = 162'b111111111101100010000000000001001011111111111101111011111111111010010010000000000001011101111111111111001110000000000011000010111111111001000000000000000001001110;
    mem[96] = 162'b111111111110010000111111111101011001111111111111001001000000000001000100111111111110110110000000000010001100000000000001011001000000000010100111111111111110010101;
    mem[97] = 162'b111111111100010110000000000000000101111111111110100100000000000001000000000000000000100011000000000001011111111111111110110010000000000000100110000000000001110101;
    mem[98] = 162'b111111111110011001111111111111001001111111111110010101111111111111011001000000000001010010111111111101010100111111111111101110000000000010001001000000000001010110;
    mem[99] = 162'b111111111101011100000000000011000000000000000000000101111111111011001110111111111010110110111111111000000101111111111111010001000000000000001000000000000001000101;
    mem[100] = 162'b111111111100100001000000000010001011000000000011011100111111111110011000111111111100101011111111111111011100000000000000111000111111111111000111000000000001010001;
    mem[101] = 162'b111111111111110100111111111111100001111111111100110110111111111111000100111111111110110001111111111101111011000000000000000000111111111100110011000000000001100101;
    mem[102] = 162'b111111111111001001111111111011100011000000000001010101000000000001011111000000000001100110111111111111100000111111111100001011000000000000001000000000000000011111;
    mem[103] = 162'b111111111101011110000000000000000001000000000000001110000000000000101100000000000000110110111111111101111011000000000001101110111111111111010001111111111111010110;
    mem[104] = 162'b111111111111111000111111111101100010111111111110110010000000000000111001000000000000110000111111111101000010000000000000001000000000000010010010111111111111101011;
    mem[105] = 162'b111111111110101000000000000010010000111111111111001100000000000000111011111111111100100101111111111111000001000000000000101000111111111101011101111111111111110100;
    mem[106] = 162'b000000000000011100111111111111110111111111111110010111111111111110111010111111111110100111111111111111011111111111111111010100000000000001011101111111111110001100;
    mem[107] = 162'b111111111111100101000000000000010010111111111110011110111111111110010110111111111111001010000000000000110011000000000001000100000000000010000101111111111111111001;
    mem[108] = 162'b111111111100100111111111111111000000111111111111000100000000000000001100111111111110001110111111111111000101111111111110111110111111111110010110000000000011011110;
    mem[109] = 162'b111111111110111101111111111111011111000000000000110001111111111110111001000000000000111011111111111100011100000000000010110000111111111100001000111111111100011101;
    mem[110] = 162'b111111111101011111111111111111011110000000000001010100111111111101101011111111111011111100000000000001011100111111111111111010111111111111100110111111111111011100;
    mem[111] = 162'b111111111101111011000000000000110000000000000011110100111111111110000110111111111101101001111111111111111000111111111101100011111111111111011110000000000001100110;
    mem[112] = 162'b000000000100111101000000001001100110000000001000000111000000001000000111000000001001011010000000000110010011000000001000110001000000000100111001000000000101000011;
    mem[113] = 162'b111111111110011011000000000001110100000000000000010100111111111101110101000000000000110010111111111110100000111111111111110010000000000001000101000000000001100110;
    mem[114] = 162'b111111111101111111000000000011110100000000000101001101000000000010101100000000000000001010000000000010001101111111111011010010111111111101110010111111111101110100;
    mem[115] = 162'b111111111111110010000000000001010000000000000000011001000000000010000001111111111101000110111111111111101011111111111110101111111111111111101011000000000010010100;
    mem[116] = 162'b000000000010000010111111111100100000000000000010011111111111111111101101000000000001000011111111111110101001111111111101111001111111111111100001111111111111000001;
    mem[117] = 162'b111111111110000110111111111110110100111111111101101111111111111101100011000000000000101100111111111010011011000000000000111100111111111110010110111111111110111011;
    mem[118] = 162'b111111111111011100111111111110100101000000000000000001000000000010101101111111111110111001111111111110101001111111111011100011111111111100111101111111111110000010;
    mem[119] = 162'b111111111110100000111111111110101000111111111110100011111111111110101111111111111111111111111111111100001100111111111111100110111111111111101000000000000000110101;
    mem[120] = 162'b000000000001100110111111111100101001111111111100111011000000000001000110000000000011010110111111111101110000111111111111011100111111111110001000000000000000111001;
    mem[121] = 162'b000000000100001100000000000011111101000000000101101110000000000100000111000000001000100100000000000100110010000000001010111011000000000100101110000000000110000100;
    mem[122] = 162'b111111111110010000111111111111011000111111111101110001111111111100110101111111111101000011000000000001001110000000000001000010111111111110111010111111111101100001;
    mem[123] = 162'b000000000000101000111111111111010110000000000000100110111111111111001101111111111011101101111111111100011111111111111101011100000000000001001110000000000000111100;
    mem[124] = 162'b000000000011001010000000000001000000000000000001000000111111111111100100111111111110011110000000000000001110111111111110010101111111111110011001111111111111010011;
    mem[125] = 162'b111111111111001111111111111110010010000000000000001110111111111101111110111111111111010100111111111111100111111111111101010100111111111101100100111111111101001110;
    mem[126] = 162'b111111111110010010111111111111000001111111111100010110000000000010101110111111111110110011111111111111100101000000000000010000111111111110111110000000000001010111;
    mem[127] = 162'b111111111011000000111111111101010011111111111110100001000000000001010111000000000000011110000000000000011010000000000001011101000000000000100001000000000000010001;
    mem[128] = 162'b000000000001101000000000000010101011111111111101010001111111111111000001111111111111100001111111111111010110111111111111101000111111111111000100000000000000110110;
    mem[129] = 162'b111111111111111111000000000000000110111111111111111010111111111111110011000000000000000010111111111111111001111111111110000000000000000000110111111111111111000011;
    mem[130] = 162'b000000000000000010000000000000000101111111111111111110111111111111101111111111111111111001111111111111111010111111111111111001111111111111111011000000000000000010;
    mem[131] = 162'b111111111111111101000000000000001010000000000000000010000000000000000110111111111111111000111111111111111111111111111111111111000000000000000011111111111111111110;
    mem[132] = 162'b000000000101000000000000000010000100000000000011101100000000000100001000000000000100001010111111111111101010111111111111110110111111111111011000000000000001100011;
    mem[133] = 162'b000000000000000000111111111111110101000000000000001100000000000000001010000000000000000101000000000000001001000000000001010100000000000011010000000000000101011010;
    mem[134] = 162'b000000000000000001000000000000001010111111111111001001111111111111111110000000000000000111000000000000001010000000000000000010000000000000000110000000000000000100;
    mem[135] = 162'b000000000001101110000000000000100011000000000000000000000000000000100000000000000010111110111111111111111000000000000000011111111111111111011110000000000000101111;
    mem[136] = 162'b000000000010011111111111111111111110000000000000111101111111111111010110111111111111110101000000000000000101111111111111011100000000000000010000000000000001101010;
    mem[137] = 162'b000000000000001010000000000000000010000000000000010001000000000000001100000000000000001111000000000000010001000000000010101000000000000010111101000000000100100011;
    mem[138] = 162'b000000000000100010111111111111110000111111111111001000111111111111111001000000000000000001000000000000000101000000000000000000000000000000000000111111111111111111;
    mem[139] = 162'b111111111111111011111111111111100010000000000000000000000000000000111100111111111111011111000000000001011000111111111111010000111111111111101001000000000000001111;
    mem[140] = 162'b111111111111111101111111111111110011111111111111111001111111111111111000111111111111111110111111111111111011111111111111111011000000000000000011000000000000001100;
    mem[141] = 162'b111111111111111011111111111111111011111111111111101100111111111111110001000000000000000000000000000000000000111111111111110100111111111111110110111111111111110000;
    mem[142] = 162'b000000000000000101000000000000000100111111111111111110111111111111110011111111111111110001111111111111110110111111111111111000111111111111110100111111111111110010;
    mem[143] = 162'b111111111111111111000000000000000100000000000000000010111111111111111110000000000000000001000000000000001001000000000000001000000000000000000100000000000000000101;
    mem[144] = 162'b000000000000000101111111111111111100000000000000000000000000000000000110000000000000000101000000000000001000000000000000001110000000000000000111000000000000000011;
    mem[145] = 162'b111111111111111110111111111111110111000000000000010011111111111111110100111111111111111010000000000000000100000000000000000110111111111111110111111111111111111110;
    mem[146] = 162'b000000000000000110111111111111111111000000000000001000000000000000000011000000000000001100111111111111111010000000000000000000000000000000000111111111111111111110;
    mem[147] = 162'b111111111111110111000000000000000110111111111111111010000000000000000010000000000000001010111111111111111011111111111111111101111111111111110010000000000000001010;
    mem[148] = 162'b111111111111111110000000000000001100000000000000000101111111111111111101111111111111111011000000000000010010000000000000001001000000000000000111000000000000001000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100111111111111111101;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule