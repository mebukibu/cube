`include "num_data.v"

module w_rom_28 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b111111111011011110111111111000011001111111111100011100111111111101001110000000000000011001000000000100000011000000000001011100000000000011101001000000000001110110;
    mem[1] = 162'b111111111011110101000000000000010101000000001000100101111111101111000110111111111011001011111111111101011001111111111000001101111111111011111111000000001000000100;
    mem[2] = 162'b000000000000010001000000000001111100111111111101000001000000000010011101000000000010101001111111111011010011000000000001000101000000000001110101111111111110001000;
    mem[3] = 162'b000000011001001001111111111111101001111111111100010001000000010101001111111111111011001111000000000001010010000000001001001101111111110001101001000000001100011101;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b000000000101001010000000000010100000111111111111111001000000000010010100111111111000010000111111111101011111111111111000010110111111110101110110000000000000000011;
    mem[33] = 162'b000000000011001000000000000000011100111111111000100101000000000100011001000000000001000011000000000000111000000000000110101011111111110100000100000000000001001001;
    mem[34] = 162'b111111111111010111111111110111100000000000000001100011000000000000110010111111111011110100000000000001110110111111111111111001111111111110000001000000000100010111;
    mem[35] = 162'b111111111110010100111111110101111000000000000110110001000000000000100110000000000000001011000000000001111001111111111110010000000000001100010100000000000111110110;
    mem[36] = 162'b111111111011001100000000000011110010000000000101110000000000000111111110111111111100010100000000000010000001000000000100111000000000000100110011000000000111110110;
    mem[37] = 162'b000000000000001010000000000000011100111111111111110110000000000011110001000000000101011110111111111110011110000000000001011111111111111101000111000000000001001100;
    mem[38] = 162'b000000000011111111000000000001011100000000000101000011111111111011001000000000000000100010000000000111110110000000000101110110000000000110101010000000001000010110;
    mem[39] = 162'b000000000010011010111111111011111011111111111010110010111111111011001111000000000100100010000000000101011011111111111000111110000000000100110010111111111101100110;
    mem[40] = 162'b000000000001010000000000000001111010000000000101011110000000001110111000111111111011111111000000000110001010000000000111110110000000000010000110000000000010101100;
    mem[41] = 162'b000000001100001111111111111110001001000000000001000000000000000000111100111111111110010000000000000010111000000000000000110010000000000011001110111111111011011001;
    mem[42] = 162'b111111110100111000000000001000101011111111111101010111000000000110000011111111111101111110000000000001101010111111111100101000000000000101100000111111111110100101;
    mem[43] = 162'b111111111110011011111111111111111011000000000010101010111111111100010100000000000011011101111111111111110101000000000100011011000000000100110001000000001101101000;
    mem[44] = 162'b111111111110011100000000000110000011111111111101001111000000000111011110111111111110011111000000000000000000111111111100001101000000000010101111000000001000011001;
    mem[45] = 162'b000000000011000001111111110101101100000000000000111001111111111111000101000000000110001100111111111000001110000000000000100000111111111100110110111111111101100101;
    mem[46] = 162'b000000000110011110111111111111001111111111111111000111111111111100100110000000000000110011000000001000001110000000000111011000000000000001001011111111111010011011;
    mem[47] = 162'b111111111111010100111111111100011111000000000110001111000000000001000000000000000010110111111111111001010100000000000001110010000000000000000110111111111110100100;
    mem[48] = 162'b000000000010100011111111111110110011000000000010101100000000000010010100111111111011110011111111110010110011111111111100000000000000000110100010111111111101110110;
    mem[49] = 162'b000000000001101111000000000110010111111111110101111111000000000100111101111111111100110000111111111101101011111111110111110110111111110110010110111111111000010001;
    mem[50] = 162'b111111111010011010000000000010100101000000000011011011000000001001110100111111111100011100111111111001110101000000000011011011111111111010111101000000000101100010;
    mem[51] = 162'b000000000001110000000000000010000101000000000110001001000000000001010100000000000110010100000000000011010101000000001000000001000000001010100000000000000101110000;
    mem[52] = 162'b111111111101110110111111111111010010000000000000001000000000001010101100000000000111101010000000000010000000000000001010000111000000000100111011000000000100001010;
    mem[53] = 162'b111111111010001100111111111101101100111111110100100000000000000100010000000000001010110011111111111101001100000000000010101110111111111110000011111111111010101000;
    mem[54] = 162'b000000000010010100000000000001000100111111111110110001000000000001110011000000000111011010111111110011110000111111111100100100111111111111011010111111110111011101;
    mem[55] = 162'b111111111010110011000000000010010101111111111111101011000000000101110100111111111010001101111111111011010100000000000001101011111111111110111110000000000011001110;
    mem[56] = 162'b111111111110110111111111111111001010111111111111000111000000000001101010000000000100011101111111111100011010000000000111010001000000000101010100000000000011011001;
    mem[57] = 162'b000000000101111110000000001101001001111111111011101110111111111011110110000000000000100010111111111010101101111111110110100111000000000010110011000000000010001011;
    mem[58] = 162'b000000000001001111111111111011101100000000001000100010111111111010001001000000000000011001000000000100010011000000001001001100000000000110011011000000000011000101;
    mem[59] = 162'b111111111101100111111111111100110010111111110110101111111111111011000001000000000100010101000000000000100111111111111100011101000000000010110101111111111101111001;
    mem[60] = 162'b111111111101101101000000000010010101111111111101001110111111111110001101000000000101110100111111110100001101111111111100100111000000000101000001111111111010100101;
    mem[61] = 162'b000000000001111010000000000101111001111111111101101010000000000010010010111111111110001111000000000101110000000000000010000011111111110011001101111111110111011010;
    mem[62] = 162'b000000000100110100000000000011101101111111111011110111111111111011000010000000000100001000111111111000110001111111111010011101111111111101111111000000000100001101;
    mem[63] = 162'b111111111110110111000000000101100101000000000000011011111111111111000011000000000001101101000000000010011010000000001000000010000000000101111010111111111010010111;
    mem[64] = 162'b111111111101010010111111111001111010000000000001111000111111111110101101111111111111001000000000000000010101000000000100111010111111111111110100111111110101111101;
    mem[65] = 162'b000000000100001000111111111111100011111111111010100100000000000001000100111111111110111011111111111101010100000000000010000101000000000001000011111111111111100010;
    mem[66] = 162'b000000000000101100000000000010111010111111111010000110000000000001101010111111111110110011111111111111010001111111111101111110000000000011100110111111111100011010;
    mem[67] = 162'b111111111010101000111111111000011010000000000010001111111111111111101011000000000110100000000000000010010001111111111011001100000000000011100111111111111100000000;
    mem[68] = 162'b000000000111000011000000001000011101000000000011001000111111111111000110111111111100101001111111111010010001111111111111011111111111111000101001111111111111001011;
    mem[69] = 162'b111111111111111001000000000000000010000000000000111101111111111010001011111111111011100011111111111110000000000000000010000100111111111011010000000000001001100000;
    mem[70] = 162'b000000000000100010111111111001000001000000000100111001111111111110101011000000000100011111111111111111001001000000000011001000111111111111101010111111111110000101;
    mem[71] = 162'b000000001000001110000000000011000100000000000001010101111111111100110100000000000001001010000000000100101001111111111111100010000000000000100100111111111101110000;
    mem[72] = 162'b000000000101010100111111111110111101000000000001000001000000000010100011111111111111000110111111111110010111000000000000001000000000000000010011111111111000111101;
    mem[73] = 162'b111111111000110101111111111011011011000000000000100011111111111110100011111111111001010100000000000100100111000000000100100110111111111011010000111111111000100100;
    mem[74] = 162'b000000000110010101000000000001010001000000000001111111111111111101100001000000000001011011111111111100101101111111111100001000000000000010010111111111111111001101;
    mem[75] = 162'b111111111111010010111111111110111001000000000100110100000000000001101100000000000001011000000000000101010110111111111101010011111111111110111010111111111010011100;
    mem[76] = 162'b000000000010001011000000000011001100000000000010111110000000000100011011000000000110001010000000000010101010000000000100111111000000000101000100000000000110011101;
    mem[77] = 162'b000000000010001001000000000100110100111111111111110001000000000011011101111111111111001011000000000001001000000000000110001001111111111011000011111111111110110101;
    mem[78] = 162'b000000000101000001000000001000100110000000000110000011000000000110101100000000000010100101000000000101101111000000000101111110000000000000001011000000000010110111;
    mem[79] = 162'b111111111111100100000000000010101100000000000011100100000000000010010000000000000011001001111111111101111100111111111110110001111111111111011000111111111100111000;
    mem[80] = 162'b111111111011000000111111111011100010000000000000111110111111111011000100000000000011011011111111111111101010000000000001100011111111111010011011111111111101111010;
    mem[81] = 162'b000000000011001101111111111101011101000000000011011000111111111110111000000000000000011110000000000100001000000000000000111111111111111011010000000000000010110101;
    mem[82] = 162'b000000000011110101000000000011100000000000000011001001000000000100100110111111111100001100000000000100110001000000000001110111111111111111101110000000000010111011;
    mem[83] = 162'b111111111111001110000000000001110101111111111101100101000000000101000100000000000001001111000000000011010000000000000110100000111111111111111111000000000100011111;
    mem[84] = 162'b111111111111000111111111111011111011111111110111110110000000000010001010111111111101010000000000000000100100111111111010101101000000000001001100000000000000100001;
    mem[85] = 162'b111111111100110100000000000101101100000000000100100001000000000010000100111111111100101100000000000011001101000000000001101001000000000001000111111111111010101001;
    mem[86] = 162'b000000000001000100000000000001111101000000000011111011000000000011101010000000000011011010000000000111000000000000001010111001000000001001010011000000001010001000;
    mem[87] = 162'b000000000011110110111111111001100111111111111010000111111111111011111000000000000000001110000000000001101011111111111100111000000000000010011011000000000000001001;
    mem[88] = 162'b111111111100111101111111110101110001111111111110100110000000000100000101111111110100111011111111110111000101111111111110111110000000000000000111111111111100101111;
    mem[89] = 162'b111111111010011101000000000011110111111111111110111110000000000000110001111111111100011010000000000010010111111111111101001000000000000001010101111111111000101110;
    mem[90] = 162'b000000000000101011000000000001100000000000000011100001000000000011111010111111111110101000111111111110001111111111111001011100111111110111100100111111111110001100;
    mem[91] = 162'b111111110110011010111111111111100110111111111001111101000000000011000001000000000001001100000000000000101100000000001011111011000000000001011011000000000100011111;
    mem[92] = 162'b111111111001111001111111111101011110111111111011000111000000000010000001000000000010001110111111111111111010111111111101110100111111111101100001111111111000001011;
    mem[93] = 162'b000000000001011100000000000000110011111111111001100111111111111111000110000000000010100111111111111111000101000000000001000110111111111101010001000000000110001011;
    mem[94] = 162'b111111111000101101111111111110001011000000000010011001000000000000111010000000000000010100111111111011110001111111111110100111000000000100011111111111111110101000;
    mem[95] = 162'b000000000000000100111111111110111110111111111110111011000000000100010001111111111011001000111111111101111110000000000000000100111111111110010111000000000011111000;
    mem[96] = 162'b111111111111110101111111111111110100111111111111110010000000000000000010111111111111111001111111111111111101111111111111101111111111111111100111111111111111110011;
    mem[97] = 162'b000000000000001010000000000000000001000000000000000000000000000000001001111111111111111011111111111111110010000000000000011001000000000000001110111111111111101111;
    mem[98] = 162'b111111111111111100111111111111101101111111111111111000000000000000001011000000000000001100000000000000000111000000000000101000000000000000100111000000000000001001;
    mem[99] = 162'b111111111111111101000000000000000011111111111111110111111111111111111001000000000000001100000000000000001000111111111111110000111111111111111101111111111111111000;
    mem[100] = 162'b000000000000000100111111111111111111000000000000000001111111111111111101111111111111111111000000000000001010000000000000001111111111111111111111000000000000000010;
    mem[101] = 162'b111111111111101111000000000000000011000000000000000001000000000000000000000000000000001001000000000000001001111111111111111001111111111111111110111111111111101010;
    mem[102] = 162'b000000000000000110111111111111111101111111111111101101111111111111111011111111111111111011111111111111110110000000000000010000111111111111111111000000000000000000;
    mem[103] = 162'b111111111111110100111111111111101101111111111111111110111111111111110101000000000000001001000000000000000110111111111111111110111111111111110111111111111111110001;
    mem[104] = 162'b111111111111100110111111111111111100000000000000000100000000000000001000000000000000000011111111111111110010111111111111111100000000000000000011111111111111111101;
    mem[105] = 162'b111111111111101110000000000000000010000000000000000100000000000000001000111111111111111110111111111111111010111111111111111110111111111111110100111111111111110000;
    mem[106] = 162'b000000000000001011000000000000001000111111111111111010000000000000000001000000000000000001111111111111101101000000000000001000000000000000001000000000000000000010;
    mem[107] = 162'b000000000000000000111111111111110111111111111111110111111111111111110000111111111111101000111111111111111111000000000000000101111111111111111111000000000000000000;
    mem[108] = 162'b111111111111111111000000000000011000000000000000000111000000000000000010000000000000010100000000000000011000000000000000011111000000000000001011000000000000001001;
    mem[109] = 162'b000000000000001011000000000000001000111111111111101010111111111111111110111111111111111010111111111111110000111111111111110000000000000000001100111111111111111100;
    mem[110] = 162'b111111111111111111000000000000001101000000000000000010111111111111110011111111111111111001111111111111101101000000000000010000000000000000010100000000000000000101;
    mem[111] = 162'b111111111111110110111111111111101110111111111111111000111111111111111101111111111111100111111111111111110000000000000000001011111111111111111101111111111111110110;
    mem[112] = 162'b000000000000110101000000000000100011000000000000011111000000000000011000111111111111110100111111111111111110111111111111100000000000000000000101000000000000011001;
    mem[113] = 162'b111111111111111011000000000000000010111111111111111000000000000000000111111111111111111010000000000000000110111111111111010100000000000000000000000000000000011010;
    mem[114] = 162'b111111111111111101111111111111101001111111111111110001111111111111110111111111111111110110000000000000001100111111111111101110111111111111111101000000000000000100;
    mem[115] = 162'b111111111111110101111111111111011111111111111111101101000000000000000110000000000000000010000000000000000111111111111111111000000000000000000110000000000000001100;
    mem[116] = 162'b000000000000001110000000000000000111000000000000011100111111111111101101111111111111101110111111111111110111111111111111110010111111111111111101000000000000100100;
    mem[117] = 162'b000000000000000010111111111111110011000000000000000000111111111111111100111111111111110010111111111111011110111111111111111100111111111111111011000000000000000010;
    mem[118] = 162'b000000000000100101000000000000010001000000000000000101000000000000001011111111111111111111111111111111111101000000000000000101000000000000001110111111111111111111;
    mem[119] = 162'b111111111111111011111111111111111110000000000000000100111111111111111100111111111111110110000000000000001001000000000000001101111111111111110001000000000000010101;
    mem[120] = 162'b111111111111101010000000000000000010000000000000001010111111111111110101000000000000000111000000000000000001000000000000100010000000000000001011000000000000000100;
    mem[121] = 162'b111111111111111011111111111111111101000000000000000100111111111111110111000000000000000000000000000000000101000000000001001010000000000000010010000000000000001010;
    mem[122] = 162'b111111111111110001111111111111111111111111111111110011111111111111101000111111111111110110000000000000000010111111111111010001000000000000001110000000000000001111;
    mem[123] = 162'b111111111111111000111111111111111100111111111111111001111111111111111100000000000000001100000000000000001101111111111111011111000000000000000010000000000000001110;
    mem[124] = 162'b000000000000001010111111111111111111000000000000001001000000000000001010000000000000001001111111111111111010000000000000010010111111111111110001000000000000001010;
    mem[125] = 162'b111111111111110010000000000000000000000000000000001101111111111111110001111111111111101001111111111111101111000000000000010100000000000000011001000000000000011000;
    mem[126] = 162'b111111111111101000000000000000000001111111111111101101111111111111111010111111111111111110111111111111110011000000000000000111000000000000000001000000000000001001;
    mem[127] = 162'b111111111111111111111111111111111111000000000000001001000000000000001000111111111111111100111111111111111000111111111111111110000000000000001000000000000000010000;
    mem[128] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[129] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[130] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[131] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[132] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[133] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[134] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[135] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[136] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[137] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[138] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[139] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[140] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[141] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[142] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[143] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[144] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[145] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[146] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[147] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[148] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule