`include "num_data.v"

module w_rom_13 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000100010001111111111111010001111111110001000100111111111010011110111111111010111111000000000010011011111111111001001110111111111111110111111111111111011110;
    mem[1] = 162'b111111010101100000000000000011010110000000001000110000111111111110011110000000000010110110000000000010000100111111010111001101000000000010011110000000000010000000;
    mem[2] = 162'b000000000001000000111111111101010111111111111111101011000000000101110100000000000010011000000000000100000110111111110111100000111111111000001000111111111110011111;
    mem[3] = 162'b000000000011011010111111101101111101000000001110110001111111111111101111000000001011011101111111111111111111111111111110001001111111101011000110000000000111111001;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b000000000000100011111111111110111100111111110110011001111111111101010011111111111011000000111111111011110011000000000001000011000000000000100000111111111110111101;
    mem[33] = 162'b000000000101101001111111110001100100000000000010100000000000000001110110000000000100000000000000000111111011111111111001000011000000000111111000111111111001101010;
    mem[34] = 162'b000000000011000000000000000000001000111111111101111100111111111011110000111111111010001110111111111011110101000000000101110111111111111010010010111111111101100111;
    mem[35] = 162'b111111111111011011111111111110011110111111110010111111000000000100011001111111111110010010000000001000111101111111111111011100000000000000111011111111111010010100;
    mem[36] = 162'b000000000010111010111111111111011011000000001100000011111111111101111011000000000010011111000000000100010001000000000110011100111111111010000110000000000101001000;
    mem[37] = 162'b111111111111110001111111110011011001111111111011001110000000000011010111000000000001011100000000000000100110111111111101011000111111111100001000111111111110101001;
    mem[38] = 162'b000000000101111100000000000100110100000000000111100110000000000010101001111111111111010110000000001001010011000000000001111101111111111110110001000000000100110100;
    mem[39] = 162'b000000000101001000111111111111111001111111111011011100000000000000011110000000000101011011000000000001111110111111111111100011111111111001010010000000000010111010;
    mem[40] = 162'b000000000000001111111111111101111101000000000110010010000000000110111000000000000100100000000000000010001110111111111111011010111111111000110010000000001001110101;
    mem[41] = 162'b111111111100101011111111111010010101111111111111110110000000000000100011111111111001101110111111111111101011000000000101100110111111111010010111000000001001001111;
    mem[42] = 162'b000000000110001100111111111101001001000000000110010101000000000001101111000000000000010101000000000011010000000000000100010001111111110111000101000000001010011010;
    mem[43] = 162'b111111111010111000111111110111010111000000001000001100000000001001011111111111111111110011111111111011011111111111111110110110111111110111110110000000000111110100;
    mem[44] = 162'b111111111110100110111111110111011001000000000101111011000000000100110000000000000111101100111111111100100000000000000011110011000000000001100010111111111101011011;
    mem[45] = 162'b111111111101110110111111111110111110000000000100011001000000000010111100000000001000011010000000000010000110000000000001100110111111111011001111111111111001001100;
    mem[46] = 162'b000000000011010000000000000001110111000000000011111010000000000010010011000000000010000001000000000001111011111111111100011110111111111110001000000000001001000100;
    mem[47] = 162'b111111110111010110000000000101001110000000000010001010111111111110001101000000000011011000111111111101010000111111111110010001111111111010111000000000000101010110;
    mem[48] = 162'b000000000101100101000000000011011100000000000000100100000000000010101010111111111010000111000000001001001010111111110110111110111111101110101010111111111001110101;
    mem[49] = 162'b000000000010000100111111110001011001111111111101001011000000000000010011000000001000100111000000000001101000000000001001001111000000000101010101111111111111101110;
    mem[50] = 162'b000000000001011000111111111001011100000000000101000001111111111110011100000000000100011110111111111101010011111111111111100011111111111110110110111111111101111111;
    mem[51] = 162'b000000000111111000000000000101010100000000000111010000000000000111000111000000000101001001000000001010100101000000000100100001000000001001010011000000001110110010;
    mem[52] = 162'b000000000011000000000000000000110010000000000010101101000000000011011000000000000001000110000000001000101011000000000110000100111111111111100000111111111111101000;
    mem[53] = 162'b111111111110111111111111111101101001000000000001111010111111111001000111111111111101000001000000000001100111000000000101000110000000000011000001000000000010110111;
    mem[54] = 162'b000000000111010011111111111100011011111111110110010111111111111111010100000000000000001110111111111101000001000000000010100000111111111011101000111111110111000110;
    mem[55] = 162'b111111110101110010111111111001010100000000000011010001111111111001111000000000000010011100111111111111100011000000000001000010000000000001010100111111111000011000;
    mem[56] = 162'b111111111010110111000000000110010101111111111101111111111111111110010111111111111010110100111111111001100010000000000111001111000000000000101010000000001001000111;
    mem[57] = 162'b000000000001111010000000000000000111000000000000001000111111111101101111111111111011000010111111111011010100000000000100100011000000000011010101111111111000000001;
    mem[58] = 162'b000000000010100010000000000001000001000000000110001100000000000100000001000000000001111100000000000001110000000000000001111000111111110111001100111111111111110101;
    mem[59] = 162'b000000000000100010000000000000000111111111111110111000000000000101000011111111111111100110111111111111000111000000000001100010000000000100011001111111111010100010;
    mem[60] = 162'b111111111000001001000000000000101011111111111010000101111111111111001011000000000110001110000000000001011111000000000101000000000000000001001101111111111100010101;
    mem[61] = 162'b000000000010011111111111111011011000000000001000100101000000000000110110000000000001111111000000000101101110000000000011101001000000000010100010000000000101110111;
    mem[62] = 162'b111111111110000010000000000100000111111111111100000100111111110100100011111111111111101111111111111111000100000000000000101010111111111011101010111111111100001010;
    mem[63] = 162'b000000000101101000000000000000100100111111111001110011111111111110110101000000000101001100000000000011101001000000000001110011000000000101001101000000000101100010;
    mem[64] = 162'b111111111101100101111111111100011001000000000011001010000000000011101010000000000001101010000000000001110101111111111101011010111111111101000100111111111101001111;
    mem[65] = 162'b111111111101010101000000000010000010111111111101010001111111111100100000000000000001011000111111111101001001000000000100011010000000000000101011000000000000001111;
    mem[66] = 162'b111111111110010001111111111010000101000000000001001101000000000011110001111111111100110100000000000010010010000000001000001101000000000011100110111111111111101001;
    mem[67] = 162'b111111111110101010000000000101110111000000000011011000000000000000111111000000000010111001000000000010101001111111110110100010000000000011011110111111111110001110;
    mem[68] = 162'b111111111010010011000000000001101000000000000001110111000000000011011000000000000010110000111111111110000100111111111100101001000000000111000100000000000010000110;
    mem[69] = 162'b111111111010111100111111111011001100000000000001101110000000000010001110000000000011011001111111111111010100000000000010010001000000000000011100111111111011001111;
    mem[70] = 162'b111111111111001100000000000010101001111111111111010100000000000011110010000000000010000111000000000101011001111111111110011000111111111011000001111111111111110000;
    mem[71] = 162'b000000000001010111000000000000010010111111111100011100000000000001010111000000000000001100111111111111110100000000000001100101111111111101110011111111111011011101;
    mem[72] = 162'b111111111000100000000000000101001011000000000000011111111111111110001110111111111111110001111111111110010100000000000000110101111111111100101001000000000111000001;
    mem[73] = 162'b111111111010101001000000000010011111111111111100100110111111111100111111111111111110110101000000000001001001000000000010100011000000000111110100111111111111011000;
    mem[74] = 162'b000000000000000011111111111111000010111111111011111100111111111110101001111111111100001000111111111111000001000000000011011011111111111110100100000000000100010111;
    mem[75] = 162'b000000000010101011000000000111001101000000001010011110000000000010101100000000001000001001000000000001010100111111111111101100111111111001101000111111111111100011;
    mem[76] = 162'b000000000000010100000000000011111100111111111110101010111111111110101001000000000100101101111111111111010000000000000101101010000000001000110011000000000101001011;
    mem[77] = 162'b000000000001000011000000000011001001111111110111011111000000000000111011000000000000111101111111111101001011111111111011001001111111111010110111000000000011101100;
    mem[78] = 162'b000000000100001100000000000011001001000000000011001011111111111110010011000000000010010011000000000001100001000000000100010010000000000010011010111111111001111010;
    mem[79] = 162'b000000000100101001111111111011001100000000000110101101000000000100011011000000000100111000111111111011101101000000000100101101111111111111110110111111111100111000;
    mem[80] = 162'b000000000011011001111111111111100001000000000001000001111111111110111000000000000011110111000000000110111011000000000010000110000000000011111000111111111111000110;
    mem[81] = 162'b000000000011100010111111111110000101000000000110100001111111111001010111000000000000001100111111111101111011111111111110101101111111111010110001000000000111101011;
    mem[82] = 162'b000000000101110001000000000111010111111111111110111000000000000001101001111111111110100101000000000100001011111111111101100010000000000000111110000000000011001001;
    mem[83] = 162'b000000000101100101000000000000011100000000000011010011000000000001110001000000000000110111000000000011010000000000000111010101000000000001001111111111111110010110;
    mem[84] = 162'b111111111000001010000000000001110010111111111111010001000000000011001011111111111100011111000000000010000110000000000110101111000000000101111100111111111100011100;
    mem[85] = 162'b111111111001011101000000000100010011111111111111100110000000000000001010000000000001110110000000000000110011000000000010100001000000000010001000111111111101101101;
    mem[86] = 162'b111111111100010001000000000010111100111111111110010101000000000001001011000000000010100100111111111111001000000000000110101111000000000110110101000000000110100010;
    mem[87] = 162'b000000000111011101111111111111011111000000000011110111000000000011000000000000000100011101111111111101101010111111111010011111000000000110001111111111110111110001;
    mem[88] = 162'b111111111111100001000000000000011101000000000001111011000000000010111010111111111001101000000000001000000001000000000000100000111111111000011001000000000100011011;
    mem[89] = 162'b111111111100111101000000000011001110000000000001100000000000000001001100000000000001100100000000000000010001111111111001101100111111111011001100000000000010000000;
    mem[90] = 162'b111111111010011101000000000011011011000000000011000010000000000001111001000000000001011001000000000001100001111111111001101110111111111111011000111111111011110111;
    mem[91] = 162'b111111110110101001000000000001000011111111111100101100000000000000111100111111111110011110111111111101100101000000000010000111000000000001011011111111111111010100;
    mem[92] = 162'b000000000000010110111111111111100111111111111101000100000000000010111111000000000010011010111111111100110100111111111000000001111111111101101101000000000010101101;
    mem[93] = 162'b111111111110100010111111111011101001111111111111101001000000000011110001000000000001110000000000000000010011111111110111111000111111111110001001111111111101110011;
    mem[94] = 162'b111111110101001111000000000101000011000000001000101100000000000011111100000000000010001000111111111011101011111111111001011010000000000000100111000000000100101011;
    mem[95] = 162'b111111111100000011000000000001111101000000000010111101111111111111100011000000000001111001111111111101110110000000000100110010000000000010010101000000000001000010;
    mem[96] = 162'b111111111111111001111111111111111010111111111111111110000000000000100011000000000000000100000000000000001111111111111111101010111111111111110110111111111111111111;
    mem[97] = 162'b000000000000001010111111111111111101000000000000000011000000000000010011000000000000011011000000000000000100000000000000010111111111111111111100000000000000001101;
    mem[98] = 162'b000000000000100001000000000000000100000000000000000000000000000000001100000000000000101010000000000000010001111111111111100110111111111111111100111111111111100111;
    mem[99] = 162'b000000000000011110000000000000010100000000000000000101111111111111110111111111111111100101111111111111110000111111111111100101111111111111101111111111111111111011;
    mem[100] = 162'b111111111111111111000000000000000100000000000000010000111111111111111100111111111111111110000000000000010110000000000000001011111111111111111001111111111111111000;
    mem[101] = 162'b000000000000000110000000000000001010111111111111110010000000000000010010000000000000000101000000000000001011000000000000100000000000000000010011000000000000000111;
    mem[102] = 162'b111111111111111000000000000000001101000000000000001110000000000000001010000000000000001001111111111111111110111111111111110100000000000000010010000000000000000011;
    mem[103] = 162'b111111111111101010111111111111110101111111111111111011000000000000010000000000000000100111000000000000001001111111111111111011000000000000001110000000000000001101;
    mem[104] = 162'b111111111111110100000000000000010001111111111111111100000000000000000010111111111111110111000000000000010010000000000000001111111111111111110111000000000000001000;
    mem[105] = 162'b000000000000000100111111111111110101000000000000001000111111111111110110111111111111110000111111111111101100000000000000001000111111111111111111111111111111111101;
    mem[106] = 162'b111111111111110101000000000000001101000000000000001100111111111111111000000000000000010100000000000000001101000000000000001001000000000000000000000000000000000101;
    mem[107] = 162'b111111111111111010000000000000000000000000000000000000000000000000000010000000000000001100000000000000000100000000000000010100000000000000001000111111111111110111;
    mem[108] = 162'b111111111111111101000000000000000101000000000000000110000000000000001001000000000000000100000000000000010110111111111111110010000000000000000010111111111111110010;
    mem[109] = 162'b000000000000100001000000000000010111000000000000000010111111111111111010000000000000000010000000000000000000000000000000001001111111111111111010000000000000000011;
    mem[110] = 162'b000000000000001011000000000000000011000000000000001001111111111111111101111111111111111111111111111111111101000000000000000101000000000000000100000000000000011100;
    mem[111] = 162'b000000000000010000000000000000000010000000000000011000000000000000011010000000000000000110000000000000000011000000000000100011000000000000011010000000000000001011;
    mem[112] = 162'b000000000000111010111111111111101010000000000001000010000000000000000100000000000000000001111111111111101110000000000000101010000000000000100010000000000000010101;
    mem[113] = 162'b000000000000000100000000000000000111111111111111110111111111111111110100000000000000000110111111111111100011000000000000001100111111111111111110000000000000000111;
    mem[114] = 162'b000000000000100011111111111111110010000000000000000111111111111111111110111111111111111110000000000000000110000000000000001011111111111111111100000000000000000000;
    mem[115] = 162'b000000000000000110000000000000000111000000000000010000000000000000001110000000000000001100000000000000011010000000000000010110000000000000001100000000000000001111;
    mem[116] = 162'b111111111111110100111111111111111110111111111111111100111111111111110111111111111111101001000000000000000100111111111111111010000000000000000010111111111111100101;
    mem[117] = 162'b111111111111111101000000000000001010111111111111111110000000000000011101000000000000001010000000000000001111000000000000000000111111111111101111111111111111110111;
    mem[118] = 162'b000000000000000011000000000000000010000000000000010001000000000000000101000000000000001010000000000000000010000000000000000011000000000000000011111111111111101110;
    mem[119] = 162'b000000000000010101000000000000001000111111111111111101111111111111111000000000000000000110000000000000000101000000000000000000111111111111110111000000000000000001;
    mem[120] = 162'b000000000000000000000000000000000001000000000000101010000000000000011101111111111111111111000000000000000110111111111111101110111111111111101101111111111111111000;
    mem[121] = 162'b000000000000000000000000000000010101111111111111110111000000000000000101000000000000001000000000000000010010000000000000000111111111111111010000000000000000011011;
    mem[122] = 162'b000000000000001110000000000000001100111111111111111010111111111111110010111111111111111111000000000000001001000000000000010101000000000000001110000000000000000101;
    mem[123] = 162'b000000000000001111111111111111110000000000000000000011000000000000001001111111111111111111111111111111111100000000000000000000111111111111111111111111111111111100;
    mem[124] = 162'b000000000000000010000000000000001101111111111111110111111111111111110011111111111111110011000000000000001010111111111111101010111111111111110001000000000000000010;
    mem[125] = 162'b111111111111110000111111111111110110111111111111101010000000000000000001000000000000001010000000000000001101111111111111110000000000000000010010000000000000001001;
    mem[126] = 162'b000000000000001110111111111111110110000000000000010011000000000000001011000000000000000100111111111111111100000000000000000010000000000000001011000000000000001100;
    mem[127] = 162'b000000000000000010000000000000000110111111111111111001000000000000000010111111111111110011111111111111110000000000000000001000000000000000001000111111111111101101;
    mem[128] = 162'b000000000000100111000000000010100110000000000011100111000000000011010100111111111111110000111111111111110000111111111111101101000000000001010111000000000000011101;
    mem[129] = 162'b111111111111111001000000000000000000000000000000000011111111111111111011000000000000001010000000000000000000111111111110111100000000000010110100000000000000001000;
    mem[130] = 162'b000000000000000110000000000000001001111111111111111111000000000000000100000000000000000010000000000000000100111111111111111101111111111111111100111111111111110101;
    mem[131] = 162'b111111111111111000000000000000000001111111111111110111111111111111111010000000000000000000111111111111111100111111111111111101000000000000000111000000000000001100;
    mem[132] = 162'b111111111111011110000000000000011100000000000000000101111111111111100101000000000000001010111111111111111011000000000000010011000000000000001000111111111111001000;
    mem[133] = 162'b111111111111110000111111111111110110000000000000001111000000000000000001000000000000000111111111111111111110000000000000010011111111111111101000111111111111111110;
    mem[134] = 162'b000000000100011011000000000101000110000000000011001010111111111111111011111111111111111111000000000000000010000000000000000001111111111111111000111111111111110011;
    mem[135] = 162'b000000000000011011111111111110001111000000000000000001000000000000000100111111111111100110000000000010010100000000000010000100000000000001001101000000000011011101;
    mem[136] = 162'b000000000000000111000000000000000010000000000000000111111111111111111111111111111111111100000000000000000101111111111111111110000000000000000111000000000000000010;
    mem[137] = 162'b111111111111111110000000000000000101000000000000001111000000000000000111000000000000000001111111111111111010000000000000000010000000000000000110000000000000000001;
    mem[138] = 162'b000000000000000101000000000000000110111111111111111110111111111111111101111111111111111011000000000000000010000000000000000100111111111111111011111111111111110110;
    mem[139] = 162'b000000000000001000111111111111111101111111111111110110000000000000000010000000000000000011000000000000000110000000000000000111111111111111111101111111111111111011;
    mem[140] = 162'b000000000010101100000000000101001011000000000101001111000000000010110001111111111101110010000000000000001100000000000000110011111111111111111100111111111101011101;
    mem[141] = 162'b000000000000000001000000000000000110000000000000000010111111111111111011000000000000000010111111111111111011000000000011110011000000000011000000000000000000110000;
    mem[142] = 162'b000000000010111110000000000101101110000000000100001100111111111111110100111111111111111100111111111111111010111111111111111011111111111111111001111111111111111000;
    mem[143] = 162'b000000000000100001000000000000010010111111111111110101111111111111111110000000000010111100000000000000001100000000000000001001000000000000101000000000000001011010;
    mem[144] = 162'b111111111111111010000000000000000011111111111111111001111111111111111111000000000000000010000000000000000011000000000000000010000000000000000100000000000000000000;
    mem[145] = 162'b000000000000000110000000000000000000000000000000001011000000000000000010000000000000001100000000000000000111000000000000000101111111111111111011000000000000000010;
    mem[146] = 162'b111111111111111011000000000000000000000000000000000010000000000000000101000000000000001000000000000000001000000000000000000100111111111111111101111111111111111111;
    mem[147] = 162'b000000000000000100000000000000001101111111111111111011000000000000000001111111111111111110000000000000000000111111111111111101000000000000001000111111111111111111;
    mem[148] = 162'b111111111111110001111111111111111010111111111111110100111111111111111011000000000000000001000000000000000100111111111111111101000000000000000101111111111111111110;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000111111111111111001111111111111110001;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule