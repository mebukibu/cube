`include "num_data.v"

module w_rom_7 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000010000111000000000100111010111111111001101000111111110110101110000000000011111010000000000011101110111111111110000000000000001000010110000000000100001010;
    mem[1] = 162'b111111111010111001000000001000001000111111110100011110000000001001011100000000000101011000000000000101001011111111111111010111111111111111111110111111111101110011;
    mem[2] = 162'b111111111111100111111111111111010001000000000000000101000000000001011001111111111000001001111111111100011010111111111110000100000000000101011000111111111111011000;
    mem[3] = 162'b000000010001100111111111111001101101000000000011101011000000000100111001111111110110001110000000001101001110000000001000101100111111111101000111000000000101000101;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111110001001001000000000100010011000000000010011001111111110000011100111111111100001001000000000000011100000000000011001001000000000101010000111111111101000111;
    mem[33] = 162'b000000000111110001111111111011110101111111111110010001000000000001010110000000000010000011111111111000110101111111111110100100000000000000000100000000000111101111;
    mem[34] = 162'b111111110101111101111111111101111101111111111000100110111111110111010111111111111100000110000000000000000010000000000110011110000000000111111011111111110111010011;
    mem[35] = 162'b000000000101011110000000000101100111000000000111000000111111110111110111000000000000010111111111111111101001111111111111010001000000000001110000111111111011101010;
    mem[36] = 162'b111111111101110100000000000100100001000000000111001101111111111100100100000000000100110010000000001010101000000000001101111111111111111011000010111111111101101100;
    mem[37] = 162'b111111111110110011000000000001011101111111111111100101000000000000100100000000000100100110000000000000000000000000001000101110111111111001110111111111111000100000;
    mem[38] = 162'b000000000111101001000000000011011111111111111110111011000000000011111001000000000001100001000000000011101100111111111111111001000000001100011001000000000000111110;
    mem[39] = 162'b000000000000001101111111111111111001000000000001000000111111111101111110111111111011011110111111111010011101111111111100110100000000000001000010000000000100000001;
    mem[40] = 162'b000000000010110111000000000000111011000000000110000110000000000001110111111111111111001001000000000111101110111111111101100011111111111111111000000000000101100110;
    mem[41] = 162'b111111111101011001111111111111100000000000000001111101000000000111010100000000000010110100000000001000100110000000000110011011000000000011100001111111110110101111;
    mem[42] = 162'b000000000011011010111111111111010100000000000000001000111111111010101001000000000001010100000000001001100111111111111001111011111111111010100000000000000000110110;
    mem[43] = 162'b000000000110001010000000000010101010000000000001000101000000000100110001000000000100010001000000000101101000000000000011110000000000000001001101111111111101010000;
    mem[44] = 162'b000000000011011101000000000100110010000000000000101011111111111011010000111111111111110000111111111101100111111111111111110111000000000011101110000000000000101111;
    mem[45] = 162'b000000000110100010000000000111111001000000000011010000111111111101001001111111111110011000111111111110101000000000000001101110111111111000010000000000000010010101;
    mem[46] = 162'b111111111100110110000000000010011100000000000000010010000000000110010100000000000010011110111111111011101111111111111010111101000000000011001010000000000100000100;
    mem[47] = 162'b111111111110011010000000000111110011111111111001000101111111111101101101000000000001100110000000000011010101000000000010001001111111111101011001000000000000100101;
    mem[48] = 162'b000000000000100010000000000001101011111111111111011110111111111100001010111111111111101011000000000100001100000000000001110100111111111100011111111111111011010001;
    mem[49] = 162'b000000000001000001111111111001100001111111111000001001111111111111010000000000000110001010000000000011001110111111111101011101111111111001100011111111111011101101;
    mem[50] = 162'b111111111001011100000000000001011100000000000001111011000000000001101101000000000000011001000000000101001000000000000001101011111111111000100110111111111000001010;
    mem[51] = 162'b000000001000100111000000000111000111000000001111011011000000000101000000000000000100010111000000000101111011000000001000001111000000000001100100000000001010001001;
    mem[52] = 162'b000000000110101010000000001000100011000000000010000011000000001000110010000000000010111101000000000100110111000000000101010100000000000011110110000000000000001101;
    mem[53] = 162'b000000000001001001000000000000011010111111111101111010111111110111110110111111111110001101000000000010010001000000000000011000111111111101101011111111111100000100;
    mem[54] = 162'b111111111000101000111111111111101110111111111101010101111111110011111000000000000001110101000000000101110011000000000100011000111111111010000100111111111011000010;
    mem[55] = 162'b000000000010100111000000000011011101000000001001011010000000000100110000111111111111010011000000000100110101111111111001010010111111110111111110111111111011000010;
    mem[56] = 162'b111111111101011011000000000001101010111111111001010110000000000001111110000000000111000011111111111011101111000000000000001001111111111111100001000000000101011010;
    mem[57] = 162'b111111110101010000000000000000000110000000000000000111000000000001001000111111111111011000000000000110010010000000000011100001111111111101011010111111111001011011;
    mem[58] = 162'b000000000111010111000000000100010011000000000101100011000000000001100010000000000100101010000000000100011000111111110110100000000000000100001100111111111011101110;
    mem[59] = 162'b111111111010000000000000000001101101000000000001100111000000000011110101111111111000100000111111110110111101000000000100011001000000000100110010111111111101010010;
    mem[60] = 162'b111111111000110000000000000110101010000000000000000110111111111000011001111111111100011001111111111100010100111111111111000010111111111111100010000000001000010101;
    mem[61] = 162'b000000000000011101111111111011100110111111111001111001000000000011010110111111111011011110000000000010001010111111111011111010000000001101110001111111111000000101;
    mem[62] = 162'b000000000100100100111111111100011101000000000101001111000000000011101010111111111100010010111111111111000011000000000101101001000000000101111001111111111101101010;
    mem[63] = 162'b111111111010101110111111111010111101000000001011100001000000001101001000111111111010101110111111111011100011000000000011111001111111111111111110000000000101000001;
    mem[64] = 162'b111111111111100111111111111011010000000000000100001100111111111000110100111111111110001010000000000110110010000000000010101000000000000010011101000000000100100010;
    mem[65] = 162'b000000000010100010111111111111011000111111111011110100000000000000100011000000000011110111000000000011110000000000000100011010111111111101110110111111111011101011;
    mem[66] = 162'b111111111111111000111111111100000001000000000101000011000000000000111110111111111001101101111111111110011000111111111111101111111111111110001100000000000011111100;
    mem[67] = 162'b111111111110101110111111111110111111000000000001111000111111111110100101000000000100100110111111111101111100111111111100111101000000000010111110000000000000011001;
    mem[68] = 162'b000000000001100001000000000001101011111111111101011110111111111110111111000000000110010101111111110111101001000000000011001100111111111001001001111111111011010000;
    mem[69] = 162'b111111111101001100111111111111100111000000000000100100111111111110001110111111111101010110111111111101011101000000000001001101111111111101110011111111111010011100;
    mem[70] = 162'b111111111110011110000000000000011011111111111111111000111111111111101101111111111110011110000000000001111101000000000001100100111111110111011011000000000100011101;
    mem[71] = 162'b000000000001001101000000000000101001111111111101100110111111111111010010111111111101111000000000000000110001000000000011000010111111111111110010000000000000101110;
    mem[72] = 162'b111111111110100111111111111100010001000000000011101011111111111000001100111111111100110100000000000000110000111111111001001110111111111011111101111111111111110010;
    mem[73] = 162'b000000000010000100111111111110111001000000000000110011111111111110011101111111111111111101111111111101011111111111111011010101111111111010101001000000000100100000;
    mem[74] = 162'b000000000010101100111111111111100100111111111100100011111111111010111100000000000011000101000000000101000101000000000000111111000000000010000101000000000001111010;
    mem[75] = 162'b000000000000000100111111111010111100000000000011001000111111111110100000111111111111101100111111111101010100000000000001010101111111111101001101000000000000011001;
    mem[76] = 162'b000000000001110001111111111111010101111111111101010100000000000100000001000000000011001110000000000100111100000000000000010111000000001010001000000000000101000000;
    mem[77] = 162'b111111111101010101111111111101111111111111111101011001111111111101011111111111111101011011111111111010010111111111111000000000000000000010010001111111111011111100;
    mem[78] = 162'b000000000100111100000000000100101100000000000010101011000000000111100110000000000110101011000000000101110110000000000010100010000000000110000110000000000011110010;
    mem[79] = 162'b111111111101111010111111111101000100111111111110000101111111111110001011111111111101011101000000000000100000111111111110000011111111111000101100111111111101111110;
    mem[80] = 162'b000000000110100010000000000001100111111111111101101111111111111111100110111111111011000110000000000100111010111111111010011010111111111111000101000000000001010101;
    mem[81] = 162'b111111111111110100000000000001001100000000000101010011111111111001011010111111111110110100111111111111111001000000000000010001111111111110000010000000000100111101;
    mem[82] = 162'b000000000001111101000000000100111001111111111010010010111111111011101011000000000100101011000000000100011110111111111101001111000000000000110000111111111101111001;
    mem[83] = 162'b000000000000011111111111111101010010000000000010100110000000000100101000000000000100110110000000000100001100000000000101110001000000000000100001000000000001100100;
    mem[84] = 162'b111111111011111111111111111100100010111111111000100010111111111101001011111111111110000110000000000000110101111111111110000010111111111001111111000000000010111011;
    mem[85] = 162'b000000000001011101000000000001010101111111111001101101111111111110100110111111111110110100111111111101100001000000000000000101111111111101111000000000000010000001;
    mem[86] = 162'b000000000000001001000000000010000011000000000001101011000000000110010001000000000110111010000000000010011000000000000110010010000000001000001001000000000111110100;
    mem[87] = 162'b111111111011101010000000000110110100000000000000011100000000000010010001111111111101100101111111110110111111000000000010011000111111111001100001111111111111111000;
    mem[88] = 162'b000000000010110110000000000001111110000000000000010100111111111011111010111111111111010101111111111101100001000000000000111101111111111111011010000000000000001000;
    mem[89] = 162'b000000000010100000111111111110101000111111111100001100000000000010101011111111111111001010000000000001101100111111111100110110111111111101110010111111111000111111;
    mem[90] = 162'b000000000010111011000000000000100011000000000111100011111111111101110100111111111100100011000000000101101101111111111101001101000000000011100110000000000001000010;
    mem[91] = 162'b000000000001110011000000000000110101111111111111101100000000000001011010000000000010110101111111111011100110000000000101001011000000000100010011000000000011101111;
    mem[92] = 162'b111111111100011101000000000110010000111111111001000110111111111110010011000000000001111000000000000001001001000000000001000100000000000001001110000000000101001010;
    mem[93] = 162'b111111111100111101111111111110110111111111111111011011111111111011010000111111111110111000111111111110010110111111111011100001111111111100101011000000000010101010;
    mem[94] = 162'b111111111101100100111111111111100101000000000001101011111111110111111001111111111011010011000000000101010100111111111101101011111111111101010001000000000010101100;
    mem[95] = 162'b000000000011011110111111111010010111000000000011001101111111111100011100111111111111100101000000000010111111111111111111101000111111111101111111000000000000000111;
    mem[96] = 162'b111111111111011110000000000000000101000000000000001100111111111111110101000000000000000100111111111111110110111111111111110001000000000000000110000000000000000111;
    mem[97] = 162'b111111111111110010111111111111101111000000000000000110111111111111110000111111111111101001000000000000000010111111111111111101000000000000000110000000000000000000;
    mem[98] = 162'b111111111111111110000000000000000000000000000000001010111111111111110111000000000000010100000000000000010111000000000000000110000000000000011000111111111111111100;
    mem[99] = 162'b000000000000001001111111111111111000000000000000010011000000000000001011000000000000000011000000000000000101111111111111111011111111111111111000000000000000000011;
    mem[100] = 162'b000000000000000100111111111111110110000000000000000110000000000000001000000000000000000000000000000000000101000000000000000001111111111111111100111111111111111111;
    mem[101] = 162'b111111111111100001111111111111101100000000000000001011111111111111111100000000000000000111111111111111111111000000000000000100111111111111110110111111111111101010;
    mem[102] = 162'b000000000000000000000000000000000110111111111111111100000000000000000000000000000000000000000000000000000010111111111111111001111111111111110100000000000000010001;
    mem[103] = 162'b111111111111110011000000000000000010000000000000000111111111111111110010000000000000000110000000000000010010111111111111100010111111111111111111000000000000001101;
    mem[104] = 162'b000000000000001010111111111111111001000000000000001110111111111111101111111111111111101010111111111111111100000000000000010100000000000000001011000000000000001010;
    mem[105] = 162'b000000000000011111000000000000001011000000000000010101000000000000010110000000000000010001111111111111111101000000000000001001000000000000000110111111111111111100;
    mem[106] = 162'b111111111111111101111111111111111100111111111111111110111111111111110101000000000000000111111111111111111100000000000000001001000000000000000100000000000000000011;
    mem[107] = 162'b111111111111110110111111111111101100111111111111101101111111111111101101111111111111110010111111111111111011000000000000011110000000000000010111000000000000010001;
    mem[108] = 162'b111111111111101010000000000000000011000000000000000010000000000000010110000000000000010111000000000000010011000000000000001110000000000000000110111111111111111101;
    mem[109] = 162'b111111111111111110000000000000000001000000000000001001000000000000000010000000000000000100000000000000001001000000000000011000000000000000010100000000000000001011;
    mem[110] = 162'b111111111111101100111111111111111100111111111111111010000000000000011101000000000000011001000000000000001100111111111111111111000000000000010100000000000000010010;
    mem[111] = 162'b111111111111100110000000000000001001111111111111111001111111111111110000111111111111110111111111111111110010111111111111101111000000000000001100111111111111110111;
    mem[112] = 162'b000000000000010101000000000000010111000000000000000101000000000000100001111111111111110010000000000000000101111111111111011001111111111111111101111111111111101101;
    mem[113] = 162'b000000000000001011000000000000000010111111111111110110000000000000001011000000000000001100000000000000000011000000000000001011000000000000001100000000000000000001;
    mem[114] = 162'b111111111111111101000000000000000111000000000000010111000000000000001011000000000000001010111111111111111000000000000000000111000000000000000010111111111111110110;
    mem[115] = 162'b111111111111110100111111111111111000000000000000000111111111111111110011111111111111111100111111111111111101111111111111100011000000000000001001000000000000000000;
    mem[116] = 162'b000000000000001111000000000000010100000000000000001001111111111111111111111111111111110010000000000000001110111111111111100101111111111111110100000000000000001010;
    mem[117] = 162'b111111111111110101000000000000000010000000000000000111111111111111110010000000000000000100111111111111111000111111111111111011000000000000010011000000000000000111;
    mem[118] = 162'b111111111111111011111111111111110001000000000000001000000000000000001011000000000000010110000000000000010001000000000000010001000000000000010011000000000000010110;
    mem[119] = 162'b111111111111101110111111111111101100111111111111110100111111111111111100111111111111110100000000000000010100000000000000001111111111111111110101000000000000000111;
    mem[120] = 162'b111111111111110111111111111111101000111111111111111101111111111111111000000000000000001010000000000000000101000000000000011001000000000000001010000000000000000010;
    mem[121] = 162'b000000000000001000111111111111111000111111111111111100111111111111101111000000000000000000000000000000001000000000000000111100000000000000001001000000000000101101;
    mem[122] = 162'b111111111111100001111111111111011111111111111111110011111111111111110001111111111111111010000000000000001110111111111111110111000000000000000001000000000000001001;
    mem[123] = 162'b111111111111111100111111111111101101111111111111100100000000000000000001111111111111111110000000000000001101000000000000000011111111111111110011111111111111111001;
    mem[124] = 162'b111111111111111010000000000000001011000000000000000000000000000000000111111111111111111110111111111111111110111111111111111111000000000000000111000000000000001100;
    mem[125] = 162'b111111111111110000111111111111111101000000000000000000111111111111111001111111111111111001111111111111111000000000000000000101000000000000011010000000000000001111;
    mem[126] = 162'b000000000000011100111111111111101100000000000000000110111111111111111110111111111111101111000000000000000110000000000000011100000000000000010110000000000000011010;
    mem[127] = 162'b111111111111110000000000000000010000111111111111101110000000000000010101000000000000001110000000000000000000111111111111111010000000000000000000111111111111110101;
    mem[128] = 162'b000000000000110100000000000000100000000000000010011011111111111111001000000000000001001010000000000000000111111111111110110101000000000000000000111111111110101011;
    mem[129] = 162'b000000000000001001000000000000001110111111111111111100111111111111111111000000000000000010000000000000000010000000000000011010111111111110101001111111111110110010;
    mem[130] = 162'b111111111111111100111111111111111110111111111111111110000000000000010000000000000000001110000000000000001001111111111111111101111111111111111001000000000000001000;
    mem[131] = 162'b000000000000011100000000000000001101000000000000001110111111111111111011111111111111110011000000000000000100000000000000000001000000000000001011000000000000001000;
    mem[132] = 162'b000000000010001110111111111111111110000000000001100100000000000100111111000000000110000000111111111111111111111111111111101111000000000000010011000000000000101000;
    mem[133] = 162'b111111111111110000111111111111111000000000000000001101111111111111111011000000000000000000111111111111111110000000000010100101000000000101100000000000000010110000;
    mem[134] = 162'b000000000000000111111111111111010111111111111111100110111111111111110010111111111111110011111111111111111110111111111111111111111111111111111101111111111111111100;
    mem[135] = 162'b111111111111010111111111111111111011111111111111011111111111111111101010000000000011110000111111111110101010000000000000110111111111111111111011000000000000000001;
    mem[136] = 162'b000000000000001000111111111111111000000000000000100100000000000000110011000000000000100001000000000000101000111111111111101001000000000000001010000000000000001000;
    mem[137] = 162'b111111111111111000111111111111111110111111111111111110111111111111110111000000000000000010000000000000000100000000000101010111000000000100000101000000000011110111;
    mem[138] = 162'b000000000000100110111111111111011000000000000000110110000000000000010000000000000000000000000000000000001100000000000000001010000000000000000011111111111111110110;
    mem[139] = 162'b000000000000111100111111111111100101111111111111110001000000000000010000000000000000110110111111111111111001111111111111011111000000000000100011000000000001100010;
    mem[140] = 162'b000000000000000100000000000000001101000000000000000010000000000000000011000000000000001101000000000000001010111111111111111001000000000000001001000000000000001101;
    mem[141] = 162'b000000000000000000111111111111111101111111111111111011111111111111110110000000000000000001000000000000000101111111111111110010000000000000001000000000000000000110;
    mem[142] = 162'b000000000000000011111111111111111111111111111111111011000000000000000001111111111111111100111111111111111110000000000000001100111111111111111001000000000000000101;
    mem[143] = 162'b000000000000000010000000000000000001111111111111111010111111111111111011111111111111111110111111111111111101111111111111111010111111111111111111000000000000000010;
    mem[144] = 162'b000000000000001001000000000000000011000000000000000010111111111111111011111111111111111100000000000000001100111111111111111101000000000000000100111111111111111110;
    mem[145] = 162'b111111111111111010000000000000000010111111111111111111000000000000000000111111111111111100111111111111111011111111111111111110000000000000010001000000000000000110;
    mem[146] = 162'b111111111111110110111111111111111111000000000000000001000000000000001010111111111111110001111111111111111010111111111111110100111111111111111101000000000000000101;
    mem[147] = 162'b111111111111111010111111111111110000111111111111110110111111111111110100000000000000000010111111111111111111111111111111111101111111111111110111111111111111111010;
    mem[148] = 162'b111111111111111011000000000000000000111111111111111111111111111111111011111111111111110100111111111111111111111111111111111111111111111111110111000000000000000000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111011000000000000000001111111111111110101;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule