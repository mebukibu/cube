`include "num_data.v"
`include "state_layer_data.v"

module add_bias_tb ();

  reg clk;
  reg rst_n;
  reg load;
  reg [3:0] cs;
  reg [12*32*`data_len - 1:0] d;
  wire valid;
  wire [12*32*`data_len - 1:0] q;

  add_bias add_bias0 (clk, rst_n, load, cs, d, valid, q);

    initial clk = 0;
  always #5 clk = ~clk;

  initial begin
    $dumpvars;
    rst_n=0; load=0; cs=`LIDLE; d={12*32{18'b00_0000_00_00_0000_0000}}; #10
    rst_n=1; #10
    cs=`LAYER0; #10
    load=1; #10
    #400
    load=0; #10
    cs=`LAYER1; #10
    load=1; #10
    #400
    $display("%h", q);
    $finish;
  end

endmodule

// layer0
// ffadbfeb6ffadbfeb6ffadbfeb6ffadbfeb6ffadbfeb6ffadbfeb6ff603fd80ff603fd80ff603fd80ff603fd80ff603fd80ff603fd80001d40075001d40075001d40075001d40075001d40075001d40075ff7f7fdfdff7f7fdfdff7f7fdfdff7f7fdfdff7f7fdfdff7f7fdfdffabffeafffabffeafffabffeafffabffeafffabffeafffabffeafffcd7ff35ffcd7ff35ffcd7ff35ffcd7ff35ffcd7ff35ffcd7ff35ffd63ff58ffd63ff58ffd63ff58ffd63ff58ffd63ff58ffd63ff580012c004b0012c004b0012c004b0012c004b0012c004b0012c004bff8f7fe3dff8f7fe3dff8f7fe3dff8f7fe3dff8f7fe3dff8f7fe3dffe8fffa3ffe8fffa3ffe8fffa3ffe8fffa3ffe8fffa3ffe8fffa3001ec007b001ec007b001ec007b001ec007b001ec007b001ec007b000b4002d000b4002d000b4002d000b4002d000b4002d000b4002dffbfffeffffbfffeffffbfffeffffbfffeffffbfffeffffbfffeffffbbffeefffbbffeefffbbffeefffbbffeefffbbffeefffbbffeefff987fe61ff987fe61ff987fe61ff987fe61ff987fe61ff987fe610029c00a70029c00a70029c00a70029c00a70029c00a70029c00a7002f400bd002f400bd002f400bd002f400bd002f400bd002f400bdffe6fff9bffe6fff9bffe6fff9bffe6fff9bffe6fff9bffe6fff9b00238008e00238008e00238008e00238008e00238008e00238008eff707fdc1ff707fdc1ff707fdc1ff707fdc1ff707fdc1ff707fdc1fff27ffc9fff27ffc9fff27ffc9fff27ffc9fff27ffc9fff27ffc9fff63ffd8fff63ffd8fff63ffd8fff63ffd8fff63ffd8fff63ffd8ffe2fff8bffe2fff8bffe2fff8bffe2fff8bffe2fff8bffe2fff8bffdabff6affdabff6affdabff6affdabff6affdabff6affdabff6a002c000b0002c000b0002c000b0002c000b0002c000b0002c000b0ffb83fee0ffb83fee0ffb83fee0ffb83fee0ffb83fee0ffb83fee0ffbe3fef8ffbe3fef8ffbe3fef8ffbe3fef8ffbe3fef8ffbe3fef8fff6bffdafff6bffdafff6bffdafff6bffdafff6bffdafff6bffdaffbb7feedffbb7feedffbb7feedffbb7feedffbb7feedffbb7feedffbbbfeeeffbbbfeeeffbbbfeeeffbbbfeeeffbbbfeeeffbbbfeee000240009000240009000240009000240009000240009000240009fff97ffe5fff97ffe5fff97ffe5fff97ffe5fff97ffe5fff97ffe5

// layer1
// ff6e7fdb9ff6e7fdb9ff6e7fdb9ff6e7fdb9ff6e7fdb9ff6e7fdb9ffa7ffe9fffa7ffe9fffa7ffe9fffa7ffe9fffa7ffe9fffa7ffe9fff893fe24ff893fe24ff893fe24ff893fe24ff893fe24ff893fe24ff6d3fdb4ff6d3fdb4ff6d3fdb4ff6d3fdb4ff6d3fdb4ff6d3fdb4ff553fd54ff553fd54ff553fd54ff553fd54ff553fd54ff553fd54ff5a7fd69ff5a7fd69ff5a7fd69ff5a7fd69ff5a7fd69ff5a7fd69ffdafff6bffdafff6bffdafff6bffdafff6bffdafff6bffdafff6bffa33fe8cffa33fe8cffa33fe8cffa33fe8cffa33fe8cffa33fe8cffa8bfea2ffa8bfea2ffa8bfea2ffa8bfea2ffa8bfea2ffa8bfea2ff3dffcf7ff3dffcf7ff3dffcf7ff3dffcf7ff3dffcf7ff3dffcf7ff4cffd33ff4cffd33ff4cffd33ff4cffd33ff4cffd33ff4cffd33ff85bfe16ff85bfe16ff85bfe16ff85bfe16ff85bfe16ff85bfe16ff40bfd02ff40bfd02ff40bfd02ff40bfd02ff40bfd02ff40bfd02ff5c7fd71ff5c7fd71ff5c7fd71ff5c7fd71ff5c7fd71ff5c7fd71ff767fdd9ff767fdd9ff767fdd9ff767fdd9ff767fdd9ff767fdd9ff733fdccff733fdccff733fdccff733fdccff733fdccff733fdccff677fd9dff677fd9dff677fd9dff677fd9dff677fd9dff677fd9dfef3ffbcffef3ffbcffef3ffbcffef3ffbcffef3ffbcffef3ffbcfff8e3fe38ff8e3fe38ff8e3fe38ff8e3fe38ff8e3fe38ff8e3fe38fee93fba4fee93fba4fee93fba4fee93fba4fee93fba4fee93fba4ff5dffd77ff5dffd77ff5dffd77ff5dffd77ff5dffd77ff5dffd77ffaa7fea9ffaa7fea9ffaa7fea9ffaa7fea9ffaa7fea9ffaa7fea9ffb2ffecbffb2ffecbffb2ffecbffb2ffecbffb2ffecbffb2ffecbffca3ff28ffca3ff28ffca3ff28ffca3ff28ffca3ff28ffca3ff28ff55ffd57ff55ffd57ff55ffd57ff55ffd57ff55ffd57ff55ffd57ff91bfe46ff91bfe46ff91bfe46ff91bfe46ff91bfe46ff91bfe46ff72bfdcaff72bfdcaff72bfdcaff72bfdcaff72bfdcaff72bfdcaffb17fec5ffb17fec5ffb17fec5ffb17fec5ffb17fec5ffb17fec5ff767fdd9ff767fdd9ff767fdd9ff767fdd9ff767fdd9ff767fdd9ff153fc54ff153fc54ff153fc54ff153fc54ff153fc54ff153fc54ff627fd89ff627fd89ff627fd89ff627fd89ff627fd89ff627fd89ff6fbfdbeff6fbfdbeff6fbfdbeff6fbfdbeff6fbfdbeff6fbfdbe
