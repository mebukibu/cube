`include "num_data.v"

module w_rom_2 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000011111000111111111111100001000000000100001100000000000101100100000000000010111000111111111110101100111111111100000000111111111101100110111111111101001101;
    mem[1] = 162'b000000000000001000111111111110100100111111110110000011111111111000101011111111111110010011111111111101111111111111110111011011000000000010101101111111111100100101;
    mem[2] = 162'b111111111111010111000000000100100011000000000000111111111111111100101001111111111110011100111111110011100101000000000010010111000000000100010101000000001000110110;
    mem[3] = 162'b111111101111100001111111001110010000111111100000000001111111110111101010111111111110110000111111101101111101000000001010111101111111110011011011111111111110110111;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b000000000011011110000000000010000100111111111101001010111111111001001000000000000100010110111111110111011101111111111110110110000000000000100011000000000100010001;
    mem[33] = 162'b000000000100100101000000000001000110111111111110000001000000000101110110000000000011010110111111111101101001000000000011101110111111111010100100111111111100110101;
    mem[34] = 162'b111111110011010100111111111111000001111111111111001111000000000100001111000000000010110100111111111101110010111111110110011101111111111111110011000000000100111100;
    mem[35] = 162'b111111110110000100111111111001011001111111111011101000111111111111111010000000000001000111111111111111010000000000001001101001000000001001011010111111111110110010;
    mem[36] = 162'b000000000001011111000000000100010011111111111101100011000000000110000010111111111010110101111111111100011110111111111101010001000000000100110000111111110111011111;
    mem[37] = 162'b000000000010110100111111111011001011111111111101110101111111111101110101000000000111010110111111111000110000000000000111011111111111111000011010111111111111001100;
    mem[38] = 162'b000000000111000001000000000011001111000000000100101011000000000101001111000000000101111010000000000000100010000000000101011010111111111100111111000000000010001010;
    mem[39] = 162'b111111111101000110000000000100000001111111111111000100000000000000010011000000000001110100111111111010110000000000000010001110111111111000110011000000001001000011;
    mem[40] = 162'b000000000011000111000000000011100101000000000000011101000000000101100111000000000000110101000000000001010010000000001100010010000000001000000000111111111101011011;
    mem[41] = 162'b000000001010001111111111110101100100111111111110111100000000000001010101111111111010010000111111111100100101000000000010000101111111111100011000000000000000011111;
    mem[42] = 162'b111111110111001000111111111001100111111111111100001001000000000011101010111111111100111000000000000001011111000000000001110011000000001000001000111111111100001101;
    mem[43] = 162'b000000000100011111000000000011111000111111111110110010000000000101100000111111111100101100000000001000010100111111111011101111111111111011111001111111111100110011;
    mem[44] = 162'b111111111001011011000000000010011111000000000001111111000000000100111000111111111110100111000000000110000101111111111111010101000000000110000010000000000100100000;
    mem[45] = 162'b000000000101111111111111111111100000000000000111011101000000000011011111111111111001100111000000000000010001111111111110001011111111111011010111000000000100110101;
    mem[46] = 162'b111111111110100101000000000100010000000000000010010001000000000110111011111111111111110101000000000100000010111111111010011110111111111100110001000000000101100111;
    mem[47] = 162'b000000000001011001000000000110110000111111111101001011000000000100000011000000000000000011000000000000100011111111111100010000000000000011101010111111111100100110;
    mem[48] = 162'b000000000010011011111111111011000110111111111111011001000000000011101001111111111100001011111111111001100100000000000000111010000000000000010110111111111110000101;
    mem[49] = 162'b111111111011100101000000001000101010000000000010011001111111110110100110000000000000111000000000000000001010111111111011001001111111111110001000000000000001010111;
    mem[50] = 162'b000000000010100101000000000001011001111111111100110111000000000000110010111111111010000001000000000111111011111111111100110101000000001010000010111111111000111011;
    mem[51] = 162'b000000001001010101000000000110110110000000000010011001000000000110111111000000001010001111000000000101100011111111111111100010000000000011000001000000000000000101;
    mem[52] = 162'b000000000101001110000000000101101111111111111111000010000000000011111001111111111111011001111111111110100001000000000011101110111111111110011101000000000011110011;
    mem[53] = 162'b000000001001000011111111111011001100111111110101010000000000000010001000111111111110010001000000000101011000111111110101001100111111111100111111000000000110010011;
    mem[54] = 162'b000000000001101001111111111100011011000000000010010011000000000001110100000000000101010100111111111100100011111111111111010001111111111110010111111111111100010110;
    mem[55] = 162'b000000000000011100111111111110011001111111111100000001111111110110111011111111111011010001111111111110011100000000000100110101000000000000001101000000000011110010;
    mem[56] = 162'b111111111111101010111111111100010010111111111011111001000000001000001000111111110101011101000000000100001000000000000101000010000000000011010001000000001001000010;
    mem[57] = 162'b000000000000011111111111111101100000111111111101100111111111111000100100000000000100101000111111111111110000000000000110101100000000000001011110000000000001011100;
    mem[58] = 162'b000000000010110101000000000000001011000000000100100111111111111111010111000000000001011100000000001000001011000000001000000011111111111000111110000000000101101110;
    mem[59] = 162'b111111110110010101000000000001100111111111111011111110111111111111000011111111111101101100000000000001111000111111111100111111000000000110001000000000000110101111;
    mem[60] = 162'b111111111001011001111111111111110111000000000011011010111111111110001101000000000110010010111111111101101111000000000010111001000000000111101110000000000000111001;
    mem[61] = 162'b000000001100111110111111111110111110111111111001010011000000000011110110111111111101000100000000001000011111111111110011000000111111111001101110111111111101101101;
    mem[62] = 162'b111111111111110001111111111110111010000000000001010111111111110111110100000000000001101101111111111110001100000000000000111001111111111110000011111111111111010010;
    mem[63] = 162'b000000000100001000111111111101110000000000000011101001111111110110110011000000000001101001000000000111101011000000000100010010000000000010110100111111111101010000;
    mem[64] = 162'b000000000000110000111111111110001111000000000000010100000000000000000101111111111101000001000000000001110001000000000000011100111111111111011111111111111111011111;
    mem[65] = 162'b000000000011111111000000000000000100000000000010110110000000000000000001111111111111001001000000000000000010000000000000000011111111111101000110111111110110010100;
    mem[66] = 162'b111111111111000101111111111111010111000000000000110000000000000011101011111111111111101110111111111011111010111111111110000111111111111110100000111111111100110010;
    mem[67] = 162'b000000000011100111111111111110010010111111111100101111111111111001011110111111111011000011111111111110001110000000000000000011000000000000100001000000000000011010;
    mem[68] = 162'b111111111001011000000000000100101001111111111110000000111111111101101111000000000000111101000000000010111101000000000010001101111111111100011111111111111111101001;
    mem[69] = 162'b111111111111101010000000000011001001111111111101010110000000000011001011000000000010110011111111111111110000111111111110111100000000000100110010000000000001001111;
    mem[70] = 162'b000000000010000110111111111111100000000000000001001010000000000000100011111111111111011000111111111101101000111111111110100101111111111100001100111111111101100011;
    mem[71] = 162'b111111111110010001000000000010111000111111111111011011000000000001110011000000000000111111111111111011011010000000000001011111000000000001001001111111111111100000;
    mem[72] = 162'b111111111111000000000000000001101110111111111100110100000000000000110000111111111111011100000000000000001001111111111010100010000000000100101101111111110111001000;
    mem[73] = 162'b000000000001101100000000000010100000111111110111011000000000000010100001111111111111000000000000000000001101000000000010000010111111111110001010111111111100111111;
    mem[74] = 162'b111111111111111010000000000000001000000000000010110010000000000010111011111111111111001100000000000010101100111111111111101000111111111100001000111111111110011001;
    mem[75] = 162'b000000000000010011111111111111011101111111111011110000000000000000001100111111111110000100111111111111001111111111111110010010111111111010101111111111111011011011;
    mem[76] = 162'b111111111111000010000000000001100000000000000001000110000000000101001111000000000011001100000000000100000100000000000110110100000000000101000110000000000010110010;
    mem[77] = 162'b111111111111100101111111111110000100111111111010100010000000000010010000000000000101000001111111111110001001111111111010001100111111111101001101000000000010011111;
    mem[78] = 162'b000000000100001000000000000100001110000000000010100100000000000110100101000000000011111010000000000010011101000000000111011011000000000011010101000000000001010111;
    mem[79] = 162'b111111111001101111000000000010011111111111111101101001000000000001010111111111111111010000000000000010001010000000000000001110111111111110111000000000000011000101;
    mem[80] = 162'b111111111101101011000000000000101111000000000001001100000000000000000100000000000000011001111111111110100000111111111110110011111111111110110001000000000000110101;
    mem[81] = 162'b111111111010010001111111111100100010000000000001110101000000000101001111000000000011000101000000000011010111111111111100010001000000000000110000000000000001001000;
    mem[82] = 162'b111111111111101011111111111111011011111111111011110100000000000001000111000000000000001010000000000010100000111111111011010011111111111100001101111111111110111001;
    mem[83] = 162'b000000000000100101000000000000101001000000000001000110000000000011110001000000000000010001111111111101100010111111111101110000111111111010100001111111111101111011;
    mem[84] = 162'b111111111101001111111111111111000111000000000000100000000000000000010001000000000000010001111111111100010101111111111000101011111111111111110111000000000010011011;
    mem[85] = 162'b111111111110010100000000000001001000000000000010000110000000000100110010000000000000101100000000000001111111111111111111010111000000000010101111000000000011001111;
    mem[86] = 162'b000000000100001110000000000011100110000000000001010111000000000001001001000000000100000000000000000010010010000000000101000001000000000001100100000000000010101111;
    mem[87] = 162'b000000000000110010111111111100110001000000000011101000111111111101110100000000000000011110111111111010001010111111111111011100111111111101011100111111111111101111;
    mem[88] = 162'b000000000001011000000000000100010100111111111000010000000000000010100010000000000010000100111111111111110011111111111111101101000000000010010100000000000011011000;
    mem[89] = 162'b111111111011000000000000000000010110000000000001101101111111111110000100000000000001011001000000000001100000111111111101111011111111111110010000111111111110100011;
    mem[90] = 162'b111111111111100001111111111001110000000000000000101000111111111110110100000000000001010110000000000011101111000000000010101101000000000001100011000000000001111001;
    mem[91] = 162'b111111111000110010111111111111100111111111111011100111111111111111110001000000000001000100000000000001101111000000000010111100000000000001000000111111111111110011;
    mem[92] = 162'b000000000001100101111111111100101011000000000010110011000000000011101001111111111101010100000000000000000010111111111100010101000000000010011100111111111100010001;
    mem[93] = 162'b000000000000010011000000000000111000111111111101011000111111111100000000111111111101011111000000000001010011000000000010100010111111111101011101000000000011000011;
    mem[94] = 162'b111111111100111010111111111111101100000000000001100100111111111110111001000000000011000111000000000000111100000000000001101110000000000001110001000000000011001010;
    mem[95] = 162'b000000000001101110111111111111001100111111111110101110000000000000100111000000000010010101111111111110001010000000000010010000111111111110011101000000000000010110;
    mem[96] = 162'b111111111111110111111111111111111110111111111111111110000000000000001001000000000000001011111111111111110010000000000000001101000000000000011110000000000000010100;
    mem[97] = 162'b111111111111111111000000000000000001000000000000000011111111111111101010111111111111110011000000000000000010000000000000001110111111111111111111000000000000000001;
    mem[98] = 162'b000000000000011010111111111111111111000000000000011111111111111111110001000000000000001101000000000000001000111111111111111011000000000000000101111111111111111101;
    mem[99] = 162'b111111111111110110000000000000000010000000000000000010000000000000001010000000000000001001111111111111110100000000000000001010111111111111111100000000000000000110;
    mem[100] = 162'b111111111111111001111111111111110111000000000000001001000000000000000110111111111111111110000000000000001110000000000000010100000000000000001100000000000000001000;
    mem[101] = 162'b000000000000001010111111111111110001111111111111101110111111111111110110000000000000000000000000000000001001000000000000000100000000000000010000111111111111110011;
    mem[102] = 162'b000000000000001011000000000000011010000000000000010111111111111111111100000000000000000100000000000000000101000000000000010010000000000000001110000000000000001001;
    mem[103] = 162'b111111111111101100111111111111110111111111111111110100000000000000000100000000000000001101000000000000001111000000000000000100000000000000001110000000000000000001;
    mem[104] = 162'b000000000000000010111111111111111111111111111111101101111111111111100111111111111111110001111111111111110100111111111111110110111111111111110010000000000000001101;
    mem[105] = 162'b000000000000010110000000000000010010000000000000000001000000000000000001111111111111111001111111111111110100111111111111101110111111111111110100111111111111110011;
    mem[106] = 162'b111111111111110110111111111111111001000000000000001010111111111111100110111111111111111101111111111111111010000000000000000100111111111111111001000000000000001000;
    mem[107] = 162'b111111111111111000111111111111101111111111111111101101000000000000000001000000000000000101111111111111111110000000000000001111111111111111111111111111111111110110;
    mem[108] = 162'b111111111111111010000000000000010100000000000000010100000000000000011001000000000000001110111111111111110011000000000000000110111111111111101101000000000000000000;
    mem[109] = 162'b000000000000000011000000000000000111000000000000000100000000000000000010000000000000001100000000000000000001000000000000000111111111111111111001000000000000001010;
    mem[110] = 162'b111111111111110101000000000000000100111111111111111001000000000000001110111111111111110100000000000000000001111111111111111101111111111111111110000000000000010011;
    mem[111] = 162'b000000000000010011111111111111111000111111111111111001000000000000010000000000000000010011000000000000000000111111111111101011000000000000001000111111111111110101;
    mem[112] = 162'b000000000000001100000000000000000101000000000000100000000000000000100000111111111111110010000000000000001101111111111111011010000000000000001110000000000000010100;
    mem[113] = 162'b111111111111110011000000000000001100000000000000000100000000000000000011111111111111111110111111111111101101000000000000001010111111111111111000000000000000011000;
    mem[114] = 162'b000000000000011010111111111111111010111111111111110111000000000000001101000000000000001100111111111111111110111111111111111111111111111111111101111111111111111000;
    mem[115] = 162'b000000000000000000111111111111111111111111111111101001111111111111101110111111111111110001000000000000001001111111111111111110111111111111111010111111111111110101;
    mem[116] = 162'b000000000000001000000000000000000101111111111111111000111111111111111010111111111111101111000000000000000001111111111111100011111111111111111100111111111111101110;
    mem[117] = 162'b111111111111101001111111111111110101000000000000001111111111111111111111000000000000001000000000000000000111000000000000001000111111111111101101111111111111101110;
    mem[118] = 162'b111111111111111011111111111111110000000000000000010111111111111111111010111111111111111111000000000000011100000000000000000110000000000000001110111111111111110101;
    mem[119] = 162'b111111111111100101111111111111111101000000000000001110111111111111110011111111111111111011000000000000000001111111111111111001111111111111111010000000000000000111;
    mem[120] = 162'b111111111111101010111111111111100111111111111111111001000000000000001000111111111111111101111111111111100101111111111111111001111111111111011101111111111111111011;
    mem[121] = 162'b111111111111110101111111111111111111111111111111110111000000000000000000000000000000000011000000000000000001000000000001101011111111111111111000000000000000010001;
    mem[122] = 162'b111111111111101101111111111111100111111111111111110000111111111111110000111111111111111111111111111111111001111111111111111111111111111111111001111111111111111110;
    mem[123] = 162'b111111111111110100111111111111101101111111111111110011000000000000000110000000000000000001000000000000000000000000000000001000111111111111110101000000000000001011;
    mem[124] = 162'b111111111111110100000000000000000011000000000000000111000000000000000000111111111111111110000000000000000001000000000000001010000000000000000110000000000000010100;
    mem[125] = 162'b111111111111110100000000000000000000000000000000000100000000000000000000000000000000000111000000000000000111111111111111111001000000000000000111111111111111111001;
    mem[126] = 162'b000000000000000001111111111111100111111111111111101101000000000000000111000000000000000100111111111111111000111111111111111000111111111111110010000000000000000000;
    mem[127] = 162'b000000000000000111000000000000010011111111111111111000000000000000010100000000000000000011000000000000010111000000000000011001000000000000100010000000000000010101;
    mem[128] = 162'b111111111111010110000000000001100101000000000001000001000000000000101110000000000000010011111111111111101111000000000000101111000000000000101011111111111110110101;
    mem[129] = 162'b111111111111110111111111111111110110111111111111110101111111111111110110111111111111110100111111111111111101111111111110111110000000000000101100000000000000011100;
    mem[130] = 162'b000000000000000001111111111111111101000000000000000010000000000000000100000000000000000110000000000000000101000000000000000101111111111111110100111111111111111000;
    mem[131] = 162'b000000000000000010000000000000000101111111111111111111111111111111111111111111111111111111000000000000000000111111111111111010111111111111111110111111111111110111;
    mem[132] = 162'b000000000010010011111111111110111101000000000001000001000000000100011110000000000010100011000000000000100000000000000000001111111111111111110111000000000000100011;
    mem[133] = 162'b111111111111111110000000000000000011000000000000001010000000000000000100000000000000000000000000000000000011000000000000001111000000000001101011000000000100001100;
    mem[134] = 162'b000000000100011101000000000000000011111111111110111011111111111111111100000000000000000010111111111111110100111111111111111010000000000000000000000000000000000100;
    mem[135] = 162'b111111111111011010111111111111010100111111111111110100111111111111011010000000000010111101000000000000100010000000000001000100111111111111011001000000000000100010;
    mem[136] = 162'b000000000000100111000000000000001100000000000010100001000000000000010000000000000010110001000000000000000010000000000001100101000000000000011010111111111111000101;
    mem[137] = 162'b111111111111111100000000000000000110111111111111110100111111111111110011111111111111110110111111111111111100000000000011000100000000000100101000000000000011110101;
    mem[138] = 162'b000000000001010110000000000001010110111111111110111000000000000000000000000000000000000001000000000000000001111111111111111101111111111111111000111111111111111110;
    mem[139] = 162'b111111111111101010000000000000101101111111111111100100000000000000101110111111111111010001111111111110111110111111111111111011111111111111101111000000000000010100;
    mem[140] = 162'b111111111111110110000000000000000110000000000000000001111111111111111100111111111111111001111111111111110110000000000000000000111111111111110110111111111111111101;
    mem[141] = 162'b111111111111111011111111111111111101000000000000000111000000000000000111000000000000000011000000000000000001111111111111111001111111111111110101111111111111110101;
    mem[142] = 162'b000000000000000010000000000000000100000000000000001001000000000000000111111111111111111110111111111111111110000000000000001000111111111111110011111111111111110001;
    mem[143] = 162'b111111111111111000111111111111111111000000000000000100111111111111110110111111111111111100111111111111111010111111111111111100111111111111111000000000000000000000;
    mem[144] = 162'b111111111111111000111111111111101111111111111111110111111111111111111001111111111111111010111111111111111000111111111111111100111111111111111101111111111111110111;
    mem[145] = 162'b000000000000000010000000000000000001000000000000000011000000000000000011000000000000000110111111111111110110000000000000000110000000000000000001111111111111110111;
    mem[146] = 162'b000000000000000001000000000000000010000000000000000011000000000000001000000000000000000101111111111111111111111111111111111111000000000000000001000000000000000011;
    mem[147] = 162'b000000000000000000111111111111111110111111111111101111111111111111111101000000000000000010000000000000000011000000000000000001111111111111111101000000000000000100;
    mem[148] = 162'b111111111111111100000000000000000001111111111111111011000000000000000100111111111111111010000000000000010001000000000000000011000000000000000010111111111111111011;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000111111111111111100;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule