`include "num_data.v"

module w_rom_24 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000101101010000000000001011110000000000000011010000000000010011110000000001010000010111111111101110001000000000010010111000000000011100110000000001011010111;
    mem[1] = 162'b111111111111110110000000001100111110111111111011100100111111111101101011000000001010111001000000000100011001000000000011101000000000001001110101111111110111000110;
    mem[2] = 162'b111111111101101010111111111100000110111111111110111110111111111100101111111111111101001110111111111111010111000000000010010011111111111011111111000000000001111001;
    mem[3] = 162'b111111111010111110000000000000011101000000000110101010111111110011010010111111101010011010000000000111010010111111110110100011000000001001100110111111111000111011;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111100000110111111101110000110111111110111011001111111111001100010111111110101011101111111111101000110000000000000001110000000000010001100000000001000000011;
    mem[33] = 162'b000000000001011100000000000010011111111111111110111000111111111101010000000000001000111111111111111101111011000000000010111010111111111011100001111111110111000011;
    mem[34] = 162'b111111110110100100111111110111101100000000000010010001111111110101011011111111110111111001111111111011010111000000000000010000111111111111111000111111111011110111;
    mem[35] = 162'b111111111100110001111111111111111000000000000101111111111111111101101000111111111110111011000000000001011011111111111011101100111111111001001101111111110101111101;
    mem[36] = 162'b111111111011010110000000000100101000000000000110000001000000000100011000000000000011100011000000000001111001111111111110000101000000000001011111000000000010000110;
    mem[37] = 162'b111111111110101110000000000000000101000000000011011000111111111100011000000000000000010000000000000011010101111111111110001111111111110111100011000000000001110101;
    mem[38] = 162'b000000000001100110000000000000010110000000000101000000000000000000010001000000000101101100000000000010000110000000000000001111000000000010010100111111111011001000;
    mem[39] = 162'b111111111001111110000000000000101100000000000100011110111111111101111000111111111101000001111111111011010110000000000010001111000000000101110110111111111111001001;
    mem[40] = 162'b000000001001110000000000000010010110000000000110011101000000000010001100000000000011000100000000000101001000111111111101101001111111111111000100000000000001011011;
    mem[41] = 162'b000000000001110111000000000000011100111111111111001011000000000000011100000000000011100100000000000101010110111111110100000100111111111110001010111111111100010100;
    mem[42] = 162'b000000000110000100111111111100110011111111111010110001000000001001001110111111111111000100111111111111001011111111111110111001000000000011100110111111111111001001;
    mem[43] = 162'b111111111110000010000000000010001111000000000101011111111111111110111011000000000110101010000000001000000011111111111110011111111111111101111001111111111110111000;
    mem[44] = 162'b111111111101110100111111110111101010000000000010000101000000000100011011000000000000001010000000000001101110000000000000001001111111111111010100111111111100100100;
    mem[45] = 162'b000000001000001110000000000001111010111111111011010010000000000001000001000000000111010111111111111101000000111111111110100110000000000011001110000000000000011100;
    mem[46] = 162'b000000000100011001111111111101100101111111111011011001000000000100101101111111111010011000111111111011110000111111111101110110000000000000111000111111110110111001;
    mem[47] = 162'b000000001000100000111111111111000101111111111101010111000000000001001100111111111111010001111111110110010000111111111110001101111111111111001010111111111001011001;
    mem[48] = 162'b111111111111100111000000000001101110111111111111010011000000000110100110000000000001011100111111111010010111111111111100001001000000000111111001000000000011010110;
    mem[49] = 162'b111111111101101100111111111111011001000000000000101010111111111011110110111111111100101101000000000011010100000000000000110000111111111111101000111111111101001001;
    mem[50] = 162'b000000000010011011000000000010100110111111111100101101111111110001100010111111111100100011000000000011100011000000000010110000111111111001111001111111111111001111;
    mem[51] = 162'b000000000011010000000000000101111001000000000110010100000000000110000011000000000110010100000000000100010000000000000110010100000000000001001001111111111101111000;
    mem[52] = 162'b000000000001010111000000000000011100000000000100110100000000000110011101000000001010101101000000001000001101111111111110111111000000000001001011111111111011100001;
    mem[53] = 162'b111111110110101111111111111111000110000000000111101011111111111100101011000000000100000001000000000000000010000000000111110111000000000000111111111111110010100000;
    mem[54] = 162'b111111111101000101000000000011100110111111111111100111000000000010000101111111111010101110111111111010110111000000000001010100000000000000000111000000000101110110;
    mem[55] = 162'b000000000010011111000000000000011011111111111100100011111111111001100010111111111001101101000000000011100011000000000000001000111111110011000011000000000000111011;
    mem[56] = 162'b111111111111111101111111111010110111000000000100011100111111111011110001111111110111001111000000000011010111111111111110010010000000000000011100000000000111110001;
    mem[57] = 162'b111111111101100100111111111110101111000000001000001100111111111001111100000000000011110111000000000000110000000000000001011010000000000001100101000000000100011111;
    mem[58] = 162'b000000000101110100111111111110001010000000000110000101000000000110101011111111111111101000000000000001110100111111111101111010111111111101101010111111110011001111;
    mem[59] = 162'b000000000111011111111111111111011000000000000010010001111111111010111101000000000000001010000000000100011110111111111010011011111111111010100001000000000001011001;
    mem[60] = 162'b000000000010011100111111111001111111111111111000101100111111111110111101000000000000110101000000000000010110000000000000001110111111110111010000111111111110011110;
    mem[61] = 162'b111111111001010000000000000100011001000000000011011100000000000010001010000000000010011100111111110110011011000000000001101111000000000000000110111111111011101000;
    mem[62] = 162'b111111111110100100111111111010101011000000000111111111000000000000000111000000000001100000000000000110000010111111111010010001111111111011110111111111110111010111;
    mem[63] = 162'b111111111101010011000000000001100010000000000001010010000000000011111110111111111110110110000000000100100100111111111100110001111111111101111000000000000100001100;
    mem[64] = 162'b111111111111100010000000000001001110111111110111000100111111111011000111111111111101011110111111111101100001000000000001111100111111111101110101000000000100110011;
    mem[65] = 162'b111111111101001110111111111100000101111111111110111001000000000001101101000000000101010010000000000000100011000000000011011010000000000010011000111111111110000111;
    mem[66] = 162'b111111111101100010111111111110100011111111111011010111000000000001101001111111111110000111111111111000111010000000000010100101111111111111001010000000000110010101;
    mem[67] = 162'b000000000100111110111111111100010101000000000001100100000000000010110101000000000001010010000000000010110110111111111110011000000000000001000101111111111101010100;
    mem[68] = 162'b111111111110011011111111111011101100111111111011111101000000000010101111000000000001011011111111111111100100111111111110111010111111111110101111000000000010100100;
    mem[69] = 162'b000000000011011011111111111010100011111111111111110110000000000000011010000000000001011001000000000001010100000000000010100100111111111010110101111111111011100110;
    mem[70] = 162'b000000000011101101000000000010101110000000000100111101111111111011011100000000000010110000000000000001110000111111111110010001111111111100111010111111111100110100;
    mem[71] = 162'b000000000010011101111111111111001001111111111111110001000000000010111110000000000001101111111111111101010011000000000010100100000000000001111100000000000001010011;
    mem[72] = 162'b111111111100010001111111111100111110000000000001101110000000000010101110111111111101011010111111111110000010111111111111111001111111111101100000111111111010110111;
    mem[73] = 162'b111111111100110010111111111110111011111111111111000011111111111110000110000000000001000111111111111011111111000000000010111100000000000010110010111111111011101101;
    mem[74] = 162'b000000000001010011111111111110001000000000000001001010000000000000111110111111111110100111111111111110111100000000000001111000111111111110101111111111111111111110;
    mem[75] = 162'b111111111101011011111111111011011001000000000001000010111111111101110110111111111110011000111111111101110011111111111010001100000000000011000001111111111100101111;
    mem[76] = 162'b000000000000000100000000000011100111111111111101010111000000000110001100000000001000011010000000000110000011000000000101010001000000000101011111111111111110001000;
    mem[77] = 162'b000000000010001101000000000011100111111111111110111011000000000011111100111111111110011100000000000100011000111111111101001011000000000011100101111111111010000110;
    mem[78] = 162'b000000000100010000000000000011111000000000000001011011000000000010110011000000000011011101000000000101101000000000000011001100000000000010111000000000000010101011;
    mem[79] = 162'b000000000011010000111111111111101001000000000101001011000000000001110001000000000001110011111111111110110101111111111011101010111111111111100100111111111100011011;
    mem[80] = 162'b000000000000110100111111111001010000111111111101111111000000000001001111111111111101100100000000000010000000000000000001000110111111111111111101111111111101011101;
    mem[81] = 162'b111111111111011001000000000010101001000000000000100010111111111011101100111111111111000101000000000010010111111111111111011010000000000000110111000000000000010011;
    mem[82] = 162'b000000000000101010111111111010101110000000000100001101000000000000001010111111111101011000000000000011010100111111111100000110111111111010011010000000000011001011;
    mem[83] = 162'b000000000011101001111111111001001010111111111111100010000000000011000101000000000010100010111111111101110001111111111101001101111111111111111100111111111101001110;
    mem[84] = 162'b000000000010100001000000000011000100111111111000010000000000000010010000000000000010111001111111111101111001111111111111100110111111111110001111111111111111010010;
    mem[85] = 162'b111111111101110011000000000100101010111111111101100001111111111110000101000000000011011101000000000001101011111111111111000010000000000010111111000000000001010110;
    mem[86] = 162'b000000000000011110000000000100011000000000000110000101000000000010100011000000000101111010000000001010100110000000000111000100000000000101101010000000000101100101;
    mem[87] = 162'b000000000000000110000000000010100001000000000100100100000000000011010100111111111110010010111111111110011000000000000000110011111111111110010010111111111010010011;
    mem[88] = 162'b111111111101111100000000000100100111111111110110110110111111111001100100111111111010101000000000000110011001111111111110011100111111110110110111111111111111111101;
    mem[89] = 162'b000000000010010000111111111100110111000000000000011011111111111110010010111111111110011001111111111100001011111111111101010100111111111101110100000000000001010011;
    mem[90] = 162'b000000000100001100111111111010001111111111111101101000111111111100111001000000000001111011000000000011010000111111111111000111000000000110101100000000000000000111;
    mem[91] = 162'b111111110111011100111111111001010011000000000001101001111111110111011000000000000010100111000000000010101111000000000101111001000000000110101010000000000100110001;
    mem[92] = 162'b111111111111000100000000000011010111000000000111001111000000000001100001000000000000000000111111111011010100111111110110010111000000000001010000111111111010101010;
    mem[93] = 162'b000000000000011110000000000011000100111111111110111010111111111110001010000000000000101000111111111100110010111111111011111101111111111111100010111111111011001100;
    mem[94] = 162'b111111111010110111000000000011001110000000000100011101111111111111111010111111111101111110111111111011010101111111111100000011111111110111001001111111111101010010;
    mem[95] = 162'b111111111111011001000000000000110100000000000001011010000000000001110110000000000000100111111111111101100010000000000100000001111111111111101100111111111110110010;
    mem[96] = 162'b000000000000000010111111111111110110111111111111110111000000000000000001000000000000000110000000000000010110111111111111111111111111111111111100000000000000000101;
    mem[97] = 162'b000000000000000011111111111111111001111111111111110111000000000000010111000000000000010000000000000000011010000000000000010011000000000000001000111111111111100011;
    mem[98] = 162'b111111111111111101000000000000000101000000000000000011111111111111111010111111111111111010111111111111111101111111111111111010111111111111111011111111111111110101;
    mem[99] = 162'b000000000000001011111111111111111110111111111111111101111111111111111000111111111111111011111111111111111001111111111111110110000000000000000011111111111111111100;
    mem[100] = 162'b000000000000001011111111111111111100111111111111111111000000000000000010000000000000001101000000000000000011000000000000000110111111111111111100111111111111111011;
    mem[101] = 162'b000000000000001111111111111111111011000000000000001010111111111111110110111111111111101100111111111111111010000000000000011100000000000000011101111111111111101110;
    mem[102] = 162'b111111111111111110111111111111111011111111111111101101000000000000000000000000000000001011111111111111111111000000000000000111111111111111111100111111111111110011;
    mem[103] = 162'b111111111111110111000000000000000010000000000000000100111111111111111000111111111111111010111111111111111011000000000000001101000000000000001011111111111111110101;
    mem[104] = 162'b000000000000000100000000000000001110000000000000000100000000000000001110111111111111111110111111111111101101111111111111111001111111111111110100111111111111111100;
    mem[105] = 162'b000000000000000110111111111111110101111111111111110110000000000000000001000000000000000001111111111111110111000000000000000111000000000000000010000000000000010001;
    mem[106] = 162'b000000000000001001111111111111110111000000000000000101111111111111110000000000000000000001111111111111111001111111111111110010000000000000000100000000000000000101;
    mem[107] = 162'b111111111111111101000000000000000100111111111111111110000000000000000001000000000000001010000000000000001101000000000000001100000000000000001110111111111111111000;
    mem[108] = 162'b000000000000001111000000000000001101111111111111111000000000000000001100111111111111111010000000000000000110000000000000100110111111111111110011000000000000001011;
    mem[109] = 162'b000000000000011000111111111111111101000000000000000010111111111111110110111111111111111001000000000000000011111111111111110100000000000000000001000000000000000110;
    mem[110] = 162'b111111111111111110111111111111111100000000000000001000000000000000000101111111111111110101000000000000010001111111111111111110111111111111111111000000000000000001;
    mem[111] = 162'b000000000000000111111111111111110011000000000000000100000000000000000001111111111111111000000000000000000111111111111111110110111111111111111100000000000000000110;
    mem[112] = 162'b000000000000101001111111111111111101000000000000110101000000000000000011111111111111111110000000000000001001000000000000000000000000000000010000000000000000100110;
    mem[113] = 162'b111111111111110001000000000000000100000000000000000110000000000000001100111111111111101100111111111111110001111111111111101110111111111111101110000000000000111010;
    mem[114] = 162'b111111111111111000000000000000000110000000000000011011111111111111111001000000000000000110000000000000001110000000000000001011000000000000000001000000000000000001;
    mem[115] = 162'b000000000000000100111111111111111000111111111111100010111111111111111100111111111111111100000000000000001010000000000000011000000000000000000000111111111111111000;
    mem[116] = 162'b000000000000001000111111111111110101000000000000000110000000000000000010111111111111111000111111111111111001000000000000000001000000000000001100000000000000001101;
    mem[117] = 162'b000000000000001011111111111111110011111111111111111000000000000000010010000000000000001000111111111111101101000000000000010001000000000000000010111111111111111110;
    mem[118] = 162'b111111111111101011111111111111111100000000000000000011111111111111111010111111111111110110000000000000001110000000000000001000000000000000000000000000000000010011;
    mem[119] = 162'b000000000000010100000000000000001100000000000000010000111111111111111100000000000000000100111111111111111111000000000000001110000000000000000010111111111111111010;
    mem[120] = 162'b000000000000001110000000000000000001111111111111101111111111111111111111000000000000000010111111111111111011111111111111111000111111111111110010111111111111111101;
    mem[121] = 162'b000000000000001100000000000000010010000000000000000001000000000000010101000000000000000001111111111111111111000000000000110101111111111111111000000000000000001010;
    mem[122] = 162'b000000000000001100000000000000010011000000000000010001000000000000001100000000000000001100111111111111110010000000000000001011111111111111111101111111111111111101;
    mem[123] = 162'b111111111111110111000000000000000110000000000000001000111111111111111111111111111111111100111111111111101110111111111111110100111111111111111100111111111111111011;
    mem[124] = 162'b000000000000001010000000000000001011000000000000000000000000000000000011000000000000000011111111111111111011000000000000001001111111111111110111000000000000001010;
    mem[125] = 162'b111111111111101001000000000000000111000000000000010000000000000000000011000000000000000100000000000000000100111111111111101111111111111111111100111111111111110101;
    mem[126] = 162'b111111111111110111000000000000000101000000000000000100111111111111111111111111111111111010000000000000001001111111111111011011111111111111100111000000000000101110;
    mem[127] = 162'b111111111111110000000000000000001000000000000000010011000000000000000000111111111111110100111111111111111101000000000000010011111111111111111011000000000000001100;
    mem[128] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[129] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[130] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[131] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[132] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[133] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[134] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[135] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[136] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[137] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[138] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[139] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[140] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[141] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[142] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[143] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[144] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[145] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[146] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[147] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[148] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule