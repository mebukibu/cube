`include "num_data.v"

module w_rom_16 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000111111000000000000011110101000000000000110000111111111100100001111111111011111011000000000000111101111111111110011100111111111001010001111111110101001001;
    mem[1] = 162'b000000000001010011000000001111011110111111110010110111111111111111100011111111111110010110000000010000000111000000000010101010111111111100000100000000001000010100;
    mem[2] = 162'b111111111101101101111111111101110000111111111111101000111111111100010111000000000000000011000000000001000011000000000011100101111111111101100101000000000001011101;
    mem[3] = 162'b000000001001111001000000010010001100000000000000001110000000001001011000111111111001110101000000001100010100000000000101101100111111111011101010000000000111010010;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111110111001000111111111101100111000000000110100100111111111000101100111111111101001111000000000010001101000000001110101001111111111011000101111111110110111000;
    mem[33] = 162'b000000000101001010111111111010111001111111111010010010000000000000110111111111111111100001000000000001101000111111111011001001000000000000110001111111111111000001;
    mem[34] = 162'b111111111110010111111111111001111011000000000000110100111111110110101111000000001000100011111111111011110110000000000000101111000000000110110010111111111111011110;
    mem[35] = 162'b111111111001010001111111111111001111000000000111101010000000000010010010000000001110110010111111110111111010000000000101111111111111110111101010111111110110100101;
    mem[36] = 162'b111111111110001111000000000010111000111111111010101001111111111110111000111111111100000100000000001000100010000000000000001101000000000000011010000000000111101000;
    mem[37] = 162'b000000000110011011111111111010011110111111111110101110111111111111000000000000000001010010000000000101001111111111111010011100111111111100010110000000001001010100;
    mem[38] = 162'b000000000001111111000000000000111001000000000011100001000000001000011111000000000100110011000000001001100010000000000000100110111111111111001111000000000110010011;
    mem[39] = 162'b000000000000111110000000000101001000000000000001011000111111111011001110000000000011101001000000000100110001000000000001100000000000000011011001111111111100101110;
    mem[40] = 162'b000000000010011100000000000011010110000000000001101110111111111111111110111111111011111010000000000010000110111111111100011111111111111111010011000000000001100010;
    mem[41] = 162'b000000000011010011111111111101110001000000000000001000111111111101100001111111111101011110000000001011010000111111111100100111000000000010111110111111111100011111;
    mem[42] = 162'b111111111110100110000000000001010000111111111110011011000000000010000110111111111100111000111111111011111011000000000101110011111111111111100110000000000111001110;
    mem[43] = 162'b111111111110110110000000000010011000000000000000011011000000000000000011000000000011010100000000001000011000111111110101011100111111111100100011000000001000010110;
    mem[44] = 162'b000000000001110101000000000001001111111111111111010110111111111101100010000000000101000111111111111110101010111111110111100101000000000000011100000000000000111111;
    mem[45] = 162'b111111111111110100000000000000000010111111111110110101000000000010101000111111111110100010000000001000101001000000000000001101111111111011100001111111111110100111;
    mem[46] = 162'b000000000010000011000000000000010000000000000010111000111111111001100011111111111110010001000000000000110100000000000000110101111111111011101000000000000000100000;
    mem[47] = 162'b000000000000110010111111111111110100000000000001000100111111110001010010000000000100111000111111110110101101000000000000110000111111111111010111111111111111101011;
    mem[48] = 162'b111111111110000010000000000010001110000000000000111111000000001001010010000000000111100110111111111011101001000000000100111001000000000011011111000000000100001011;
    mem[49] = 162'b000000000010011000111111111010100110111111111000000001111111111110100100111111111110110111000000000101101101111111111011100101000000000101010110111111111100111110;
    mem[50] = 162'b000000000010001010111111111110100001000000000010010000000000000010001011111111111111000110111111111011111011000000000011110001111111111100100000000000000010010011;
    mem[51] = 162'b000000000110001010000000000101011101000000000101000010000000000101001101000000000111000100000000000111110100000000000001111001000000000111011101000000000010100010;
    mem[52] = 162'b000000000110010011111111111111010000000000000011100111000000000100110010000000000010001000000000000010001000000000000101010010000000000001111111000000000011011101;
    mem[53] = 162'b000000000001000010000000000011011101111111111011101100111111111010001111000000000101010100000000000100011010000000000001101000111111111000110001111111111111011101;
    mem[54] = 162'b000000000110001000111111110111111111111111111101011111000000000011111111111111111110000000111111111110011110000000010000101111000000000000011110111111111110001110;
    mem[55] = 162'b111111111111000111000000000000110100000000000101110001000000000100100111000000000001101001111111111111111000000000000010110111111111110110011101111111111101100100;
    mem[56] = 162'b000000000001011110111111111101101101000000000110100111111111111110110001000000000000100001000000000000101011111111111111010011111111110111011100111111111100111000;
    mem[57] = 162'b000000001010111010111111111001111001111111111101101010000000000100001001000000000100111110111111111100100001111111111100100111000000001100011001111111110110001101;
    mem[58] = 162'b000000000011000101000000000000001110000000000100101111000000001000110110000000000000110011000000000011001010111111111101110101111111111011110100000000000101010110;
    mem[59] = 162'b111111111010111110000000001010000011111111110111000110000000001001100000111111111110111100000000000001010110000000000001000110000000000001010100111111111010010011;
    mem[60] = 162'b111111111101111101111111111010010011000000000001100010000000000001100111111111111110111110111111111001111000000000000011101000111111111110101111111111111000011011;
    mem[61] = 162'b000000000000011100000000000000001111111111111011111101111111111001111111111111111100001010000000000011111101000000000011000110000000000111010101000000000001100110;
    mem[62] = 162'b111111111011110010000000001000101001000000000001100001111111111000101011000000001000111111111111110101001100000000000100100110111111111111100111111111111110100001;
    mem[63] = 162'b111111111000010100000000000110001101000000000000011000000000000010011100000000000101010011000000000010000011000000000000011000111111111110010101000000000011000000;
    mem[64] = 162'b000000000011010101000000000001100010000000001000100100000000000000110101000000000000010100000000000111111001000000000110000101000000001000100010000000001000001011;
    mem[65] = 162'b000000000010110110000000000010001101000000000101101001000000000011110101000000000010100100000000000101100001000000000100011111000000000010101011000000000111101011;
    mem[66] = 162'b000000000100011100111111111110001111000000000100001100000000000010000110000000000001100101000000001000000101000000000100101111000000000111111001000000000110000011;
    mem[67] = 162'b000000000001100111000000000010101001000000000010001001111111111101011001000000000010100011000000000110000100000000000111111011000000000110100001000000000100101011;
    mem[68] = 162'b000000000001110010111111111111101010000000000001000010000000000010001000111111111111001111111111111111010011000000000001100011000000000011101111111111111111101100;
    mem[69] = 162'b000000000001001000000000000100011010000000000101111100000000000011110100000000000110001011000000000000110110000000000000011101000000000100011010000000000010011111;
    mem[70] = 162'b000000000011001001111111111110100010000000000100001100000000000001100101111111111111100000000000000100001001000000000110001111000000000010011100000000000011011101;
    mem[71] = 162'b000000000111010110000000000011010011000000000011011000000000000001111111000000000110010000000000000111110111000000000111011000000000000111000010000000001010010100;
    mem[72] = 162'b000000000101011010000000000010111101000000000111110101000000000001100010111111111101110111000000000001100010000000000011101101000000000000001111000000000010110101;
    mem[73] = 162'b000000000010100110111111111001111001111111111100101110111111111100111001111111111101101011000000000001110011000000000101100011111111111110000010000000000010001011;
    mem[74] = 162'b000000000000001010000000000001010000000000001000110111111111111111101000000000000100110101000000000010000000000000000010110010000000000010101001000000000101010011;
    mem[75] = 162'b000000000010011011000000001010110000000000010000111001000000000011110111000000000110011010000000000010100010000000001010001001000000000100001101000000000110011100;
    mem[76] = 162'b000000000111011101000000001000011010000000001110011001000000001000110111000000001100011011000000001101011001000000001100011010000000010000000111000000010001011101;
    mem[77] = 162'b000000000010000101000000000110110010000000000110101000000000000100111000111111111111001000000000000111101101000000000000011001000000000111011001000000000100101001;
    mem[78] = 162'b000000001100000010000000001011110101000000001101001111000000001000110110000000001000111110000000001111101010000000001111100101000000001010010100000000001110101100;
    mem[79] = 162'b000000001000010101000000000100011111000000001001011100000000000010001011000000000100001101000000000111010111000000000111101100000000001000111011000000001001011001;
    mem[80] = 162'b000000000010111101000000000011000100000000000111000000000000000000001101111111111111110101000000000010101110000000000010010101000000000000011001000000000110011111;
    mem[81] = 162'b000000000001111111000000000001000011000000000011010111000000000001000100000000000001101110000000000110001000000000000010100000000000000101001110000000000111001111;
    mem[82] = 162'b000000000010000011000000000001011110000000000110001001000000000011100101000000000010101010000000001010001101000000000100100101000000000010001010000000000100000101;
    mem[83] = 162'b000000000101101011000000000110011110000000010000000000000000000010110110000000000011000100000000000111100011000000001000101111000000000100110111000000000101100001;
    mem[84] = 162'b111111111101111101000000000001010101000000001000100011111111111110000000000000000000010001000000000010110011000000000110001110000000000100110010000000000100100101;
    mem[85] = 162'b000000000100110111000000000101111000000000000110111011000000000100100101000000000001111000000000001010100100000000000011111101000000000111010100000000000100101101;
    mem[86] = 162'b000000000111100011000000001011001111000000010010110100000000001010001110000000001111010110000000010011000101000000010100010011000000010110000001000000011000010110;
    mem[87] = 162'b000000000010001011111111111101101100000000000001101010111111111110111110111111111100111011000000000000010010000000000110011100000000000010111010000000000101001011;
    mem[88] = 162'b000000000000100111000000000011100001000000001001011010000000000011000101000000000001101110000000000011111101111111111111000010000000000000000111000000000101010001;
    mem[89] = 162'b000000000001110101000000000000110011000000001010101110111111111111110100000000000001100111000000000011011001000000000100111011000000000001101101000000000101111101;
    mem[90] = 162'b000000000111110101000000001001000010000000001101001001000000000100011010000000000100011010000000001001001010000000000100111110000000000111110111000000001011111011;
    mem[91] = 162'b000000000011100100000000000101100111000000001011001100000000000100101111000000000110010001000000001000000100000000001011010000000000001010110010000000001101011010;
    mem[92] = 162'b000000000010011001000000000001011001000000000100111110000000000011011001000000000011111010000000000110000000000000000110000001000000000110100010000000000011100000;
    mem[93] = 162'b000000000000101100111111111111000010000000001001100010111111111110110000111111111101100001000000000011010111000000000001100010000000000100110010000000000010000011;
    mem[94] = 162'b000000000010111100000000000000011110000000000010110010000000000011010010111111111110000011000000000001111111000000000010000010000000000011100101000000000110001001;
    mem[95] = 162'b000000000000111011000000000011101101000000001000010111000000001000010000000000000011010111000000000100101101000000001000011110000000001001010101000000000101100001;
    mem[96] = 162'b000000000010101111000000000001010011111111111010011010111111111101001000000000000001001011111111111001100010000000000001000001000000000000100010111111111110011000;
    mem[97] = 162'b000000000001011110111111111110011011000000000010111111111111111110001101000000000000010001000000000010110100111111111111101011000000000010110010111111111111110001;
    mem[98] = 162'b111111111111010111111111111101011110000000000001000101000000000001000011111111111110100100111111111111011111000000000000101010000000000001000011111111111111101110;
    mem[99] = 162'b111111111111000001111111111101101001000000000000001101111111111010000011000000000000011001000000000001101100111111111011001111000000000000011010000000000000001100;
    mem[100] = 162'b000000000110101100000000000010100111000000000110010110111111111111100110000000000010000101000000000001001001111111111110011100111111111111110000000000000001111011;
    mem[101] = 162'b000000000010011001111111111111011010000000000001111100111111111100100111111111111100110101000000000000110100111111111100111111000000000001100001000000000001101101;
    mem[102] = 162'b111111111101111010000000000000001001111111111111110101111111111100010000111111111110110010111111111100101110111111111111000101111111111110111010000000000101011101;
    mem[103] = 162'b000000000001010101111111111111011101111111111110111000000000000001000110000000000001011110111111111100110101000000000000110010111111111001011010111111111111100110;
    mem[104] = 162'b111111111101111111111111111111111101111111111111010100000000000000010010111111111111110001000000000001011100111111111110111111111111111111010100000000000101011111;
    mem[105] = 162'b111111111010111110111111111101100011000000000000010000111111111111010001111111111101100100000000000010001111111111111101011111111111111111110111111111111110000110;
    mem[106] = 162'b111111111100101001111111111110000000000000000011100001000000000001101010111111111101111100111111111111000011111111111110010101111111111011010101111111111011100000;
    mem[107] = 162'b111111111111000000111111111010100100111111111100110101111111111101111010000000000010000101000000000000010010000000000010010001111111111110100100000000000010000110;
    mem[108] = 162'b111111111100111001000000000000000001000000000001101100000000000000000100111111111110100000000000000001101000111111111101011100111111111111011100111111111111110011;
    mem[109] = 162'b000000000000100101111111111110110001111111111100111000111111111110000001111111111110010000111111111111001100111111111111110011000000000000101110111111111101111011;
    mem[110] = 162'b000000000100110001111111111101011001000000000000010100000000000010000011000000000000000001111111111111101101000000000000011111000000000001100100000000000010100010;
    mem[111] = 162'b000000000001100110111111111110011111000000000000111010111111111111011110111111111011100001000000000001101111000000000001001101000000000000010110111111111110001100;
    mem[112] = 162'b000000001010011100000000001011010100000000001101111001000000001000101000000000001000110000000000000101101010000000001000010001000000001001111010000000001101011000;
    mem[113] = 162'b111111111100100100000000000010011110000000000001011010111111111011110110111111111111100000111111111110010010111111111111111111111111111101000111000000000000111111;
    mem[114] = 162'b000000000011101100000000000000110110000000000000110100111111111111001001000000000000111010111111111110000110111111111111111000111111110100010110111111110110110001;
    mem[115] = 162'b000000000011011010000000000010010101000000000000101111111111111011001011111111111110110000111111111110011111111111111111101000111111111111110011000000000001100000;
    mem[116] = 162'b111111111110011101111111111111111000000000000010011111000000000000111100000000000001000011000000000000000110111111111111100100000000000100110101111111111111001001;
    mem[117] = 162'b111111111111101101111111111110101110000000000101111001000000000001100111111111111101010010111111111100010000111111111111001100000000000000001001000000000100100010;
    mem[118] = 162'b111111111110111100111111111110110011111111111101001100111111111100111010111111111111100100111111111011110100111111111111001010111111111110110011111111111110111100;
    mem[119] = 162'b111111111101000110111111111110000100111111111110100100111111111111011011111111111111101111000000000001101011111111111111000110111111111110001011111111111101001000;
    mem[120] = 162'b000000000001111111000000000000011111000000000011001010111111111111111111111111111011111111000000000001110100000000000000111011111111111111000101111111111111000001;
    mem[121] = 162'b000000001001011000000000001000000000000000000110101100000000000111101001000000000100001111000000000111010110000000001000010001000000001010111111000000010011010001;
    mem[122] = 162'b111111111011000110111111111111100111111111111100010001111111111101110110000000000010100011000000000000010001000000000010011010111111111111111000111111111011000011;
    mem[123] = 162'b000000000000100010000000000001000100111111111011100101111111111000010001111111111110100011111111111101100110111111111110100011000000000010110000111111111101000110;
    mem[124] = 162'b111111111111000010000000000010011000111111111101101000111111111111000010000000000000000010111111111101110111000000000001011011000000000000000100111111111100010110;
    mem[125] = 162'b111111111001101000000000000001000001111111111101110010111111111101111110111111111000111111111111111101100011111111111110101110000000000001100100111111111101010100;
    mem[126] = 162'b111111111111111010111111111110100000000000000000100101111111111110110110111111111011111111000000000000000110111111111111111100111111111110000011000000000000000100;
    mem[127] = 162'b000000000000101011111111111011100010000000000000000010111111111101000101111111111110010111111111111010101010000000000000101110111111111111010101111111111101111010;
    mem[128] = 162'b111111111111111101000000000010010001000000000101101000000000000100100010000000000001001111000000000000001111111111111111110111000000000000100010000000000000101101;
    mem[129] = 162'b111111111111101111111111111111101110111111111111110110000000000000001001111111111111110011000000000000000001000000000000011110111111111111100001111111111111101111;
    mem[130] = 162'b111111111111110100111111111111110011111111111111110001111111111111110111000000000000001110000000000000000110000000000000001110111111111111110101111111111111111100;
    mem[131] = 162'b111111111111111110111111111111110000111111111111110111000000000000000000111111111111101001111111111111101101111111111111101100111111111111100110111111111111111011;
    mem[132] = 162'b000000000000010000111111111111100101000000000000001110000000000000001001000000000000001110111111111111110110000000000000010101000000000000000010111111111111011001;
    mem[133] = 162'b111111111111101111111111111111101101000000000000000101000000000000001011111111111111111111111111111111111100000000000000011010111111111110111001111111111111111110;
    mem[134] = 162'b000000000010011110000000000010110111000000000101011010111111111111111110000000000000000110111111111111110100000000000000000000111111111111111110000000000000000110;
    mem[135] = 162'b000000000000010110111111111111110110000000000000011001111111111111110101000000000000000110000000000010001111000000000000001000000000000000010011000000000100111100;
    mem[136] = 162'b000000000000000000111111111111111100000000000000000100000000000000000110000000000000001000000000000000000101000000000000011001000000000000001101000000000000001001;
    mem[137] = 162'b111111111111110001111111111111111001111111111111110101111111111111110100111111111111111100111111111111101000000000000000000101000000000000001010111111111111111100;
    mem[138] = 162'b111111111111111110111111111111101110000000000000001000000000000000000100111111111111111010111111111111110011111111111111111000111111111111100010111111111111110111;
    mem[139] = 162'b111111111111111100000000000000001011000000000000001011000000000000000101111111111111111111111111111111110101000000000000000000000000000000000000111111111111111111;
    mem[140] = 162'b000000000011100101000000000100111000000000000100010010000000000011001010111111111111100101000000000001010001111111111111110010000000000000010111111111111101101011;
    mem[141] = 162'b111111111111101011111111111111110110000000000000000001111111111111110111111111111111110110111111111111110000000000000101001110111111111111111000000000000010111100;
    mem[142] = 162'b000000000011100110000000000101011001000000000100011111111111111111101001111111111111100110111111111111100111111111111111111001111111111111111001111111111111111001;
    mem[143] = 162'b111111111110111110000000000000101000000000000000001110000000000000101101000000000001100111111111111111110001000000000000100001111111111111111001000000000001100010;
    mem[144] = 162'b111111111111101011111111111111110101111111111111111111111111111111110101111111111111101111000000000000000001111111111111111111000000000000000001111111111111101011;
    mem[145] = 162'b000000000000000101111111111111111111111111111111111110000000000000010010111111111111111110111111111111111100111111111111101000111111111111111011111111111111101101;
    mem[146] = 162'b000000000000000000111111111111111010111111111111111000000000000000001100000000000000010000000000000000001110000000000000000100000000000000001011000000000000001110;
    mem[147] = 162'b000000000000000110000000000000000000111111111111111010000000000000000101000000000000000010000000000000001011000000000000001010000000000000000101000000000000000010;
    mem[148] = 162'b111111111111110011111111111111110111111111111111110001111111111111101001111111111111101011111111111111111101111111111111101101111111111111110110111111111111101110;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111010111111111111110101111111111111101111;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule