`include "num_data.v"

module w_rom_26 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000110000100111111111110110100000000000001000110111111111111000010111111111111011011000000000100000110000000000110001110000000000100111100111111111100011010;
    mem[1] = 162'b111111011001001000000000000000101011000000000000001000111111111110011101000000001010011111000000000010010111111111000100111011111111110100000111111111111111011001;
    mem[2] = 162'b000000000100010101111111111111111101111111111100001111000000000000001001111111111010010101111111111111000010111111111110100110000000000010001100111111111100110000;
    mem[3] = 162'b111111100001011001111111010111010100111111110110011101111111011010111000111111101001110100000000000100000100111111001001101101111111100011111000111111110110110101;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111100000000111111111101111011000000000110000011000000000011101110111111111111001111111111110101110001000000000001001101111111111011101000000000000110101110;
    mem[33] = 162'b111111111001111010111111111011010010000000000001000011000000000100100010000000000011111111000000000000000100000000000001011100111111110110010111111111111101110101;
    mem[34] = 162'b111111111100011110111111111110101110111111111110101011111111111011000011000000000000000101000000000100010001111111111011001000111111111010101100000000000101010000;
    mem[35] = 162'b111111111111001110111111111101101011111111111010100110111111110001000011111111111010111001111111111010111100000000001001001010000000000000010110111111111001111001;
    mem[36] = 162'b000000000010001001000000000000101111000000000001110100000000000111011110000000000101011100000000001010100010111111111101010101111111111111010101111111110010101000;
    mem[37] = 162'b000000000111010000000000000011001010111111111100110001111111111101001000000000000001010000000000000011111011111111111011011001000000000001011101111111110110001010;
    mem[38] = 162'b000000000001001110000000000011100111000000001010000111000000000001111110000000000110101110111111111110110101000000001010001110000000000100111100000000000000110010;
    mem[39] = 162'b000000000100010101000000000010010101111111111101111110000000001000010001111111111010010011000000000001001000000000000011101101111111111101001111000000000000011001;
    mem[40] = 162'b000000000110110110000000000011011110000000000100100011000000001000110000000000000001111001000000000010010001111111111011100101111111111110111011111111111101110110;
    mem[41] = 162'b000000000110111100000000000100110101000000000001010001000000000000110000111111111101010000111111111101111101000000000001110101111111111010011110111111111011110100;
    mem[42] = 162'b000000000011101000000000000000000101111111111011001011111111111100110111000000000111111100111111111011110000000000000000000011000000000001110011111111111110001000;
    mem[43] = 162'b000000000110001101000000000110100101000000000111011010111111111100010111000000000111000100000000000100110011111111111011100110111111111110000100111111111111101001;
    mem[44] = 162'b000000000001100000111111111011011101111111111101100000000000000001101110111111111010010101000000000011000111111111111101100101111111111110101100111111111110111000;
    mem[45] = 162'b000000000100111010000000000011101011111111111111101010111111111101000011000000000101100010111111111001010110000000000110010110000000000001110101111111111001001001;
    mem[46] = 162'b000000000000011010111111111110101110000000000100001010000000000010111111000000000101001001111111111110100100000000000110000011111111111100110100111111111010000111;
    mem[47] = 162'b000000000001000001111111111001011011000000000010010100000000000010011100000000000000000100000000000001100101111111111110001010000000000001011000111111111010110011;
    mem[48] = 162'b111111111100100111111111111001010011000000000110111110111111111101011010000000000010001101111111111000001101000000001001111111111111111110011001111111111110000101;
    mem[49] = 162'b000000001101101000000000000100101000000000000101010110111111111011011000111111111111100001000000000001100110000000000010101001111111110011100001111111110010000100;
    mem[50] = 162'b000000000100110010000000000001101110000000000111011100111111111010011111111111111001011011111111111000011100000000000100111010000000000001000101111111111110010000;
    mem[51] = 162'b000000000110110110000000000011011100000000000110011001000000001011001010000000000010111010000000000110000111000000000110010010000000001000101010111111111101101110;
    mem[52] = 162'b000000000011100101000000000011000110111111111101011001000000000100011101000000001010000000000000000011100100000000000110011011000000000100111101000000000001010000;
    mem[53] = 162'b111111111111100100000000000000011100111111110111001110000000000010110010000000000101111111000000000001001110111111111100001111111111111100010011000000001010100011;
    mem[54] = 162'b111111111111111101000000000100100110111111111110111100111111111100101010000000000001111111111111110001110111000000000000100000000000000001100111000000000101111011;
    mem[55] = 162'b000000000011100010000000000111111001000000000101011010111111111100010000111111111010001010111111111110111100111111111101011011000000000001001000111111111100101110;
    mem[56] = 162'b111111111100111111111111111111110101111111111001110010000000000000001000000000000000000110111111111100101000000000000010111000000000000111100110000000000000011100;
    mem[57] = 162'b111111111011101111000000000000110110000000000100000000111111111011111111111111111101001001111111111111000011000000001101110000111111111011110110000000000001111100;
    mem[58] = 162'b000000000010100011000000000110110001000000000001111000111111111111101111000000000001001110111111111010101100000000000001100111000000000100101101111111110110101010;
    mem[59] = 162'b111111111101101001111111111101111101111111111101101011000000000100110001111111111101101111000000000111100110111111111011110100000000000110101010111111110110001111;
    mem[60] = 162'b111111111111111011111111111001010110111111111011000101111111111000000000111111111111101011000000000001101111111111111001000111111111111011011010000000000000000111;
    mem[61] = 162'b111111111101111000000000000110011110000000000000000011000000000001100110111111111110100000111111111110100001111111111101010011111111110111111010000000000111000100;
    mem[62] = 162'b000000000110110001000000001010100110111111111110000000111111111110011100111111111100100010111111111000011011000000000001100101111111111111000011000000000011101100;
    mem[63] = 162'b000000000110011000000000000001011110111111111111000000111111111110111100000000000100110010111111111011001100111111111010111011000000000001111110111111111101000100;
    mem[64] = 162'b000000000100111110111111111101100101111111111101100111000000000011000011111111111111110011111111111110110110111111111011000101000000000100001111111111111110000100;
    mem[65] = 162'b000000000011001111000000000011111111000000000000000010000000000001100001000000000011011010111111111011101001000000000000000011000000000000110000000000000110110101;
    mem[66] = 162'b000000000001010110111111111100101010000000000001001010111111111100011001000000000001000010111111111110110110111111111110101100000000000001000101000000000000011011;
    mem[67] = 162'b111111111111010010000000000101001001111111111001101101000000000010101101000000000010111000111111111010100110000000000000000001111111111000100011111111111001010000;
    mem[68] = 162'b000000000010101110000000000000100100111111111111100011111111111110001001111111111011011010000000000000100100000000000001110110000000000010111001000000000010101010;
    mem[69] = 162'b000000000100001011000000000101010001111111111101100000111111111100001101000000000100000100111111111101001110111111111110001000111111111101001001000000000000110110;
    mem[70] = 162'b000000000001000011000000000000010001111111111100101000000000000011010111000000000101101000000000000000111000000000000010000100111111111111011001111111111101011101;
    mem[71] = 162'b000000000010100011111111111110001100111111111111100000111111111111001100000000000011101000000000000101111001000000000011101110000000000100011010111111111110101011;
    mem[72] = 162'b000000000001010101000000000000000011000000000010011001111111111101111100000000000001011011111111111011100001111111110111011100000000000001001110000000000100111001;
    mem[73] = 162'b111111111111100010111111111111011111000000000101111110000000000001001111111111111101001100000000000101100101000000000011001000000000000001000101000000000010111001;
    mem[74] = 162'b000000000101100101111111111101001111111111111111001111000000000011101010111111111011100010000000000000011010111111111001111000000000000010011010111111111100001110;
    mem[75] = 162'b000000000110110100000000000001101010111111111111111100111111111100001000111111111110101110000000000110100111111111111001100111111111111111001100111111111110010011;
    mem[76] = 162'b000000000000000101000000000100001010000000000001010001111111111111100100111111111110000101000000000010011000000000000001100100111111111110000100000000000001010100;
    mem[77] = 162'b000000000000101111000000000000110110000000000000101011111111111111100101000000000010101110000000000010010011000000000001101000111111111000110001000000000001010000;
    mem[78] = 162'b000000000010011101000000000010110011000000000011101000000000000101001011000000000010010000000000000100010100000000000110000010000000000110000111000000000100101100;
    mem[79] = 162'b000000000011010110111111111101110111000000000000011000111111111011011110111111111111101011000000000101001111111111111010111101000000000000110100111111111011001010;
    mem[80] = 162'b111111111110010000111111111110110100000000000010110110000000000010101111000000000110001000000000000110010110000000000001111010111111111001111111000000000000001100;
    mem[81] = 162'b000000000010010001111111111101001001111111111010110100000000000001101010000000000001111010000000000011001110111111111100000000000000000011110110000000000000000011;
    mem[82] = 162'b000000000100011111111111111101011011000000000000000011111111111111101111000000000011101110111111111100100110111111111100001110000000000101001111111111111011000000;
    mem[83] = 162'b111111111001111010000000000000011101111111111111001001111111111101001101111111111100110010111111111100110011111111111110110100000000000011010000000000000011010101;
    mem[84] = 162'b111111111110000100111111111001100001000000000011110000000000000001000111000000000000110000111111111101000110111111111011001001111111111111101100111111110110110010;
    mem[85] = 162'b000000000010110111000000000001111111000000000100001100000000000011110011111111111110000101000000000011111101000000000101111010111111111011000110000000000110110011;
    mem[86] = 162'b000000000000010011000000000011111001000000000111110100111111111111010100000000000100100101000000001000011010000000000100010001000000000100010111000000000101011111;
    mem[87] = 162'b000000000000001100111111111101100111000000000000010011111111111111000011000000000001001011111111111101101100111111111100100011000000000001111000111111111110101110;
    mem[88] = 162'b111111111011000011111111111100000010000000000001011101111111111110001110000000000001110000111111111100011001111111111001000010000000000100101110000000000100000010;
    mem[89] = 162'b000000000010110010111111111100001011000000000001101110000000000000010001000000000000100111111111111110111111000000000001111110000000000011000110111111111110110010;
    mem[90] = 162'b111111111011001010000000000001101101000000000100110110111111111111111011000000000000001101000000000001111101000000000001110110000000000000101100000000000010101110;
    mem[91] = 162'b000000000011110101111111111111101101000000000000100110000000000001011111000000000100011100000000000000010000000000000011001010000000000010001100000000000001010011;
    mem[92] = 162'b111111111111010010111111111110000011111111111111010000000000000011010000000000000000100100000000000000111110000000000010001000111111110101010111000000000000010000;
    mem[93] = 162'b000000000011101100111111111000111110111111111110110010111111111001001110000000000000010010111111111111001010111111111100110000000000000101111000000000000001001010;
    mem[94] = 162'b111111111111010100000000000010011111111111111110110100000000000101010010111111111111101111000000000011101100000000000000000110000000000010011101000000000010101111;
    mem[95] = 162'b111111111111010001000000000000010100000000000010010100111111111111000010111111111101111100000000000010010010111111111111011100111111111001101110000000000000001000;
    mem[96] = 162'b000000000000001000111111111111111111111111111111110101111111111111110100111111111111110101000000000000000011000000000000000100111111111111110110111111111111110100;
    mem[97] = 162'b111111111111111000000000000000000001000000000000000101111111111111111101111111111111110101111111111111101100000000000000001101000000000000000100000000000000000101;
    mem[98] = 162'b000000000000001000111111111111111101000000000000000100111111111111110111000000000000000001000000000000000011111111111111111101000000000000010010000000000000001101;
    mem[99] = 162'b000000000000001100111111111111110111000000000000001110111111111111111000111111111111111111111111111111111000111111111111111011000000000000000100111111111111110001;
    mem[100] = 162'b111111111111111000000000000000000110000000000000000001000000000000001010000000000000000011000000000000001011000000000000001000111111111111111101111111111111110010;
    mem[101] = 162'b111111111111110011111111111111110110111111111111111110000000000000000111000000000000001000000000000000001011111111111111101101111111111111110011000000000000001001;
    mem[102] = 162'b111111111111111000000000000000000110111111111111110010111111111111110110111111111111101101111111111111101000111111111111111010000000000000000000111111111111111011;
    mem[103] = 162'b111111111111111110111111111111110100111111111111101100111111111111011010111111111111111011000000000000010010111111111111101101000000000000000110111111111111111011;
    mem[104] = 162'b111111111111111001000000000000010101000000000000001111000000000000000100111111111111110110111111111111111000111111111111111100111111111111101111111111111111111000;
    mem[105] = 162'b000000000000001111111111111111110111111111111111111011000000000000000110111111111111101101111111111111110110000000000000000101111111111111110000111111111111011000;
    mem[106] = 162'b000000000000000001000000000000001100111111111111111001111111111111101111111111111111101010111111111111101011111111111111100110111111111111110000111111111111101110;
    mem[107] = 162'b111111111111111100111111111111110110111111111111111010111111111111101011111111111111110110111111111111101101111111111111110101000000000000100001000000000000010001;
    mem[108] = 162'b111111111111111111000000000000000111000000000000000001000000000000000110111111111111111011111111111111111101111111111111111101111111111111110100111111111111110010;
    mem[109] = 162'b111111111111111011000000000000000100111111111111111100000000000000001100111111111111111011111111111111111101111111111111111011000000000000000100000000000000000100;
    mem[110] = 162'b111111111111110100111111111111110010111111111111110101000000000000000010000000000000000110111111111111111110000000000000011001000000000000000001000000000000001110;
    mem[111] = 162'b111111111111101100111111111111110001111111111111110110111111111111110100000000000000001000111111111111110100111111111111111011000000000000010000000000000000010100;
    mem[112] = 162'b000000000000000000000000000000001111000000000000011011000000000000011111111111111111111000000000000000011110000000000001000011111111111111111100000000000000000101;
    mem[113] = 162'b000000000000011001111111111111111111111111111111110110000000000000000000000000000000000101000000000000000110111111111111111001111111111111110111000000000000001001;
    mem[114] = 162'b000000000000000100111111111111111101000000000000001101000000000000001001111111111111111001111111111111111110000000000000000011000000000000000010000000000000000100;
    mem[115] = 162'b111111111111101110111111111111111000111111111111101101111111111111101001000000000000000001111111111111110000000000000000001001000000000000001011000000000000011000;
    mem[116] = 162'b111111111111111000000000000000001010000000000000011110111111111111101010111111111111101110111111111111111000111111111111110011111111111111111010111111111111110001;
    mem[117] = 162'b111111111111111010000000000000001001000000000000000011111111111111011001111111111111110010111111111111101101000000000000001000000000000000010000000000000000000011;
    mem[118] = 162'b000000000000001110111111111111101111111111111111111010000000000000011001111111111111111010111111111111111010111111111111110100111111111111110001111111111111111100;
    mem[119] = 162'b111111111111111010000000000000000011111111111111111100111111111111111111111111111111101101111111111111111100111111111111101010111111111111110101000000000000000010;
    mem[120] = 162'b111111111111101100111111111111110001111111111111110111111111111111110110111111111111101001000000000000001100000000000000010010000000000000010001000000000000000111;
    mem[121] = 162'b000000000000000111111111111111110101000000000000010010111111111111110011111111111111111010000000000000001011111111111111000000000000000000010010000000000000001001;
    mem[122] = 162'b111111111111111101000000000000000101000000000000000001111111111111110000111111111111110000111111111111110110111111111111101100111111111111110011000000000000001110;
    mem[123] = 162'b111111111111111110000000000000000000000000000000001111111111111111111101000000000000000001000000000000000101111111111111110000111111111111111111111111111111111000;
    mem[124] = 162'b111111111111111010111111111111111011000000000000000011000000000000000111111111111111111100000000000000000100111111111111111101000000000000000000111111111111110110;
    mem[125] = 162'b111111111111101110111111111111111010000000000000000000111111111111011010111111111111101110111111111111100111000000000000000011000000000000010011000000000000011000;
    mem[126] = 162'b111111111111111011111111111111110110111111111111111010111111111111111111111111111111101100111111111111011111111111111111111110111111111111111001111111111111111011;
    mem[127] = 162'b000000000000001101000000000000000110000000000000001010000000000000001011111111111111111111111111111111110010000000000000000010000000000000000011111111111111111100;
    mem[128] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[129] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[130] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[131] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[132] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[133] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[134] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[135] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[136] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[137] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[138] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[139] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[140] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[141] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[142] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[143] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[144] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[145] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[146] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[147] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[148] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule