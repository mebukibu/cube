`include "num_data.v"

module w_rom_19 #(
    parameter filename = "../data/data162/weight162_0.txt",
    parameter integer dwidth = 9*`data_len,
    parameter integer awidth = 8,          // 2^8 = 256 > 5*32 = 160
    parameter integer words = 5*32
  ) (
    input wire clk,
    input wire [awidth - 1:0] addr,
    output reg [dwidth - 1:0] q
  );

  (* ram_style = "block" *)
  reg [dwidth - 1:0] mem [0:words - 1];

  always @(posedge clk) begin
    q <= mem[addr];
  end

  initial begin
    //$readmemb(filename, mem);
    mem[0] = 162'b000000000011000100111111110011111110111111110111101111111111110110011000111111111000101110000000000011101101000000000000100010111111111111100010111111111001100001;
    mem[1] = 162'b111111101101010001000000000110010001000000000111001001000000000010010111000000000100110011111111110100011111111111111010001110000000000101010000000000000010000100;
    mem[2] = 162'b111111111101101001111111111100110101111111111101010011111111111100110110111111111100011011111111100001010000111111111001010100111111101011100101111111111000110011;
    mem[3] = 162'b111111111101010110111111011001111101111111111010101110111111110101011011000000000101110010000000000100110010111111110111011111111111110100100000000000000011101110;
    mem[4] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[5] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[6] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[7] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[8] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[9] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[10] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[11] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[12] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[13] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[14] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[15] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[16] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[17] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[18] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[19] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[20] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[21] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[22] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[23] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[24] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[25] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[26] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[27] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[28] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[29] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[30] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[31] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[32] = 162'b111111111011001111111111110100011010111111111011001101000000000111110101000000000001000101000000000010000100000000001001111010111111111100000010111111110101110010;
    mem[33] = 162'b000000000110000010000000000111100010111111101110101000111111111011110111000000000100000111111111110110110001111111111110011100000000000101101000111111111100100100;
    mem[34] = 162'b111111110111101011111111111000110010000000000000001110000000000110010100111111111101000001000000000000011111111111111101011101111111111101011100111111111100000111;
    mem[35] = 162'b111111111100110110000000000001011000000000000000011110111111110010001111111111111110111101111111111011100010111111111110010000111111111100010100000000000001000110;
    mem[36] = 162'b000000000101111111000000000000110110000000000001010101000000000001100001111111111011110101000000001000101001111111111110001010000000000100010010000000000111100100;
    mem[37] = 162'b000000000010000111000000000101001100111111111011110110000000000010000101111111111010101111000000000000110001000000000010110010000000000001000100111111111000011111;
    mem[38] = 162'b000000000100100001000000000010101001000000000010001110000000000101000001000000000110000000000000000011011101000000000011001001000000000001000000111111111110100110;
    mem[39] = 162'b111111111111111010111111111101001011111111111011110001000000000011101111111111111100111010000000000101100101000000000101100000111111110111001010000000001001001100;
    mem[40] = 162'b000000000100111001111111111111100010000000000101000100000000000010100111000000001000000001000000000101001011000000001011010000000000000000111101000000000011111001;
    mem[41] = 162'b111111111110011110111111111101111000111111111101000111000000000100111111000000000010000001000000000111000000000000000011000011000000000101011011111111111110000100;
    mem[42] = 162'b000000000011110010111111111100001110000000001001000010000000000101101100000000000100010101000000000000000101111111111000100110000000000100011011000000000110100111;
    mem[43] = 162'b111111111101000110111111111101000101000000000101100011111111111100001010000000000111111011000000001000001011000000000010110011000000000001101110111111111111101000;
    mem[44] = 162'b111111111100110010111111111100110010000000000001100011111111111011111110111111111110000100111111111001011001000000001001010111111111111101010111000000000000100101;
    mem[45] = 162'b000000000100100100111111111011111000111111111100101011111111110111111000111111111111111010000000000011100111000000000100000101000000000101011101000000000111001011;
    mem[46] = 162'b111111111011000000000000000000111101111111110110111101111111111101100011000000000110110000111111111111101001000000000110010111111111110101111110000000000111111011;
    mem[47] = 162'b111111110111101110000000000010011100000000000001001111000000000110001101000000000011000010111111111110100001111111111110010101111111111010101100000000000010100110;
    mem[48] = 162'b111111111110110100000000000001011110000000001000101100111111111101110010000000000010001100000000000001001100000000000010001101000000000001101001000000000000001110;
    mem[49] = 162'b000000000100101000111111111011100011000000000011110010111111110010010101000000000010010111000000000001010111111111111101011010000000000101000000000000000000111011;
    mem[50] = 162'b111111111110111000111111111010011111000000000010111111111111111010111001000000000100111011000000000010101111000000000100001000000000000100000110000000000110000000;
    mem[51] = 162'b000000000011100111000000000100111001000000000001011100000000001001000001000000001010010100000000000011110011000000000111001011000000001110111100000000010010110010;
    mem[52] = 162'b111111111100111101000000000100000001111111111111101100000000000111011111000000000001110101000000001000101100000000000001100101000000000111000010000000001010010101;
    mem[53] = 162'b111111111101001100000000001001010110111111111011101110000000000011001100000000000000011101111111110110010100111111111100011111000000000001110101000000000010001110;
    mem[54] = 162'b000000000001100100111111111110000010111111111011110000000000000011010000111111111110001001000000000000010011000000001010101101000000001011001010111111111010010101;
    mem[55] = 162'b111111111100000011111111110011010010000000000101110011000000000001010000000000000110000101000000000000110001111111111000111101000000000010001111111111111010101110;
    mem[56] = 162'b111111111010101101111111111100100101111111111110000111111111111011100010111111111010010100111111111100000000000000000000101111000000000011101000111111111111011110;
    mem[57] = 162'b111111111101111111000000000111111001111111111100100100000000000101010010000000000011011111111111110101001110111111111000111101000000000010101100111111111110000111;
    mem[58] = 162'b111111111101011111111111111111100110111111111100010111000000000100011111000000000101100101000000000010000111111111111111110010000000000001010111000000000000001100;
    mem[59] = 162'b000000000010010011000000000001100101000000000101110111000000000011000001111111110101100111111111111010010110111111101111110001111111111110001001111111111101100110;
    mem[60] = 162'b111111111111100100111111111111010101000000000001001101111111111100100010111111111010100010000000001000001100111111111010110011000000000000010011000000000100110101;
    mem[61] = 162'b111111111111111001000000000000100111111111111101110110000000001000100101000000000000000101111111111110011000111111111100000011000000000011110100000000000001111111;
    mem[62] = 162'b111111111111100111000000000010001110000000000001110110000000000001000011111111111111010010111111111010100111111111111101010101111111111010111001111111111001011001;
    mem[63] = 162'b000000000110011110000000000111000100111111111111000100000000000000111110000000001100010011111111111011100010000000001001001111000000000101100001000000000001000111;
    mem[64] = 162'b111111111101111011111111111001010011000000000110010110000000000010101011000000000011001001000000000001000010111111111110000011000000000011100000000000000100000100;
    mem[65] = 162'b000000000001110011111111111110111111111111111100110000111111111110101000000000000100001100111111111001111101000000000100000010000000000010011000111111111011110000;
    mem[66] = 162'b111111111001101000000000000011000001000000000000010111111111111101010110000000000001110010111111111001000011111111111111101110111111111110011101111111111110110111;
    mem[67] = 162'b111111111010100001111111111110111101111111111100110011111111111100100011111111111101110010000000000011111011111111110101110110111111111111100110000000000010000000;
    mem[68] = 162'b111111111111000001000000000101100001111111111110011110111111111100001111111111111101011000111111111101101101000000000001111100000000000001010111111111111010010100;
    mem[69] = 162'b111111111101101011000000000011010111000000000101101101111111111110111000000000000101110111000000000100100011111111111110101011111111111101111000000000000001101111;
    mem[70] = 162'b000000000000100100000000000010111110000000000101000101000000000001100110000000000100111011000000000010101001111111111100100100000000000011010110111111111110011100;
    mem[71] = 162'b111111111010110001000000000010011010111111111011000101000000000011100111111111111110011111000000000010100001000000000101000100111111111000001010111111111111011110;
    mem[72] = 162'b000000000011111010111111111111001000111111110110111111000000000110100000111111111110010001111111111001100101111111111001101001111111111101111011111111111100100010;
    mem[73] = 162'b111111111010110001111111111110110010000000000010100110000000000001101101000000000101011110111111111110001001111111111010100010000000000001000010111111111111101001;
    mem[74] = 162'b111111111101000010111111111101010110111111111110111101111111111010011011111111111011001111111111111010010010000000000000110011111111111101010110111111110110000101;
    mem[75] = 162'b111111111100011010000000000001100110000000000010001001000000000111110010000000000000010011000000000001110001000000000101001110111111111100111001000000000101110111;
    mem[76] = 162'b000000000100010101111111111110100110000000000101101100000000001001010001000000000100001101000000000000001111000000000010100101000000000111101000000000000100100010;
    mem[77] = 162'b000000000000101111111111111000100101111111111010110100111111111110010110000000000001010001000000000000100111111111111011001011000000000001010100000000000001010001;
    mem[78] = 162'b000000000010001010000000001001001001000000000111011000000000000101111101000000000011011111000000000111011000000000001011001111111111111110111001111111111001010011;
    mem[79] = 162'b000000000111000001111111111100010110000000000100111111000000000111100110000000000010010011000000001000000010111111111011001101000000000011011110111111111000001100;
    mem[80] = 162'b000000000110100010111111111001110111000000000000100011000000000010100010000000000011100110111111111110101001000000000000010110111111111110011011000000000001101111;
    mem[81] = 162'b000000000101110011111111111101110000111111111011010111111111111000111110111111111110001001000000000100000010000000001000101111111111111101101010111111110110100100;
    mem[82] = 162'b111111111111010000000000000100000001000000000100010010000000000001000100111111111100110011111111111110101001111111110111011111000000000100000100111111111011000101;
    mem[83] = 162'b111111111110001000000000000110101110000000000100010111000000000010001010111111111110001111000000001000111010111111111111100001111111111100000001000000001000111110;
    mem[84] = 162'b000000000000000100111111111100001001111111110100001001000000000000011011111111111111101110111111110111111001111111111110111100111111111111011111000000000001101100;
    mem[85] = 162'b111111111111010100000000000111111011111111111111100010111111111101111100111111111101011001111111111111000110000000000011101000000000000001010011000000000101011100;
    mem[86] = 162'b111111111111110011000000000001011100000000000011100001000000000011010011000000000110000100000000000110101100000000001011001101000000000011001100000000000100110100;
    mem[87] = 162'b111111111111011001000000000000001101111111111100100011000000000010110111111111111111100010111111111111001001111111111110101011111111111110111010111111111101110110;
    mem[88] = 162'b111111111000011001111111111111010101111111111001001000000000000001101011111111111101101101000000000000001111000000000011100101111111111000101100111111111111010011;
    mem[89] = 162'b000000000110011110111111111100010011111111111100001011000000000010110100000000000000010000111111111011101111111111111111101010111111111001001010000000000101010110;
    mem[90] = 162'b111111111101110111000000000001100011111111111010001000111111111100100011000000000010110101000000000001010000111111111110011010000000000001110101000000000001010100;
    mem[91] = 162'b111111111011110111000000000011000101000000000011010010000000000011110000000000000101110100111111111111001100111111111101000110000000000011100011111111111111010000;
    mem[92] = 162'b000000000000001001000000000100111010111111111100111110111111111100010101111111110101101000000000000101011110000000000100011110000000000010010010111111111111011011;
    mem[93] = 162'b000000000000000011000000000000110000111111111101011111000000000000101000111111111111011011111111111100101111000000000000100000111111111011001011111111111101011100;
    mem[94] = 162'b111111111011011000111111111101010101000000000010010111000000000001111111000000000101010000000000000110111011000000000110110010111111111010110110111111111001100001;
    mem[95] = 162'b111111111010101010000000000001111110111111111110110010000000000011010110111111111101111111000000000010100111000000000111100011000000000001001000111111111111010000;
    mem[96] = 162'b111111111100110111111111111110011010000000000001001010000000000011100010111111111101110000000000000010010111111111111101110011111111111101111110111111111101111111;
    mem[97] = 162'b000000000001001100000000000000110110111111111111000011000000000000110110000000000010000010111111111100110011000000000001000100111111111111011111111111111011100000;
    mem[98] = 162'b111111111100100001111111111111101000111111111111010001111111111101011111000000000000101100111111111111000100111111111110111110000000000010110011000000000000111001;
    mem[99] = 162'b111111111101111000111111111111001101000000000000000111111111111110010010000000000000111100111111111111011011000000000001010101111111111110000000000000000010101001;
    mem[100] = 162'b000000000001001001000000000001010100000000000000110111000000000010111011111111111101110100000000000010110101111111111111011101111111111111101000000000000001110001;
    mem[101] = 162'b111111111111110011111111111101010010111111111111001110000000000001001110000000000000001110000000000001101000111111111011010100111111111100010011111111111110010111;
    mem[102] = 162'b111111111010010010111111111110100110000000000000000010111111111111100111000000000000010111111111111100110101000000000000000000000000000001000111111111111111001000;
    mem[103] = 162'b111111111111101001000000000001011110111111111111000101111111111111111011000000000100001111111111111101101101111111111110101100000000000000101101000000000011001010;
    mem[104] = 162'b000000000010111110000000000010101111000000000001101100111111111100000001000000000010101001000000000000011000000000000000010111000000000000000010111111111101101110;
    mem[105] = 162'b111111111111010100111111111101010110111111111111001010111111111110110011111111111111011011111111111101011111000000000000001010111111111100110110111111111100101000;
    mem[106] = 162'b000000000010111001111111111110110000000000000000110110111111111111001100111111111110001110111111111100110011111111111110001101111111111110111001111111111100100100;
    mem[107] = 162'b111111111111000110111111111111011000000000000000101100111111111111110001111111111110010110000000000001000000111111111100100001000000000001011011111111111110100111;
    mem[108] = 162'b111111111111001011000000000000101001111111111111001101000000000100110100000000000000101011000000000010011110111111111101011111000000000001001100111111111101111010;
    mem[109] = 162'b111111111110110001111111111110000100111111111010100011111111111110111111111111111110001000111111111111101010111111111101010000000000000000011110000000000000011010;
    mem[110] = 162'b111111111111100011111111111101101101000000000000001111111111111101110100111111111110100101111111111110001011111111111100011110000000000000011100111111111110100000;
    mem[111] = 162'b111111111110111001111111111011101110000000000000000000111111111100101110111111111111111101000000000001110111000000000000100011111111111111011111000000000010110010;
    mem[112] = 162'b000000000110010110000000000101100101000000000100100001000000001001100100000000000101100111000000000111011001000000001011111100000000000111001100000000000001111000;
    mem[113] = 162'b111111111111010100111111111110011101000000000011111111111111111111000010111111111111110000000000000100001000000000000001101011111111111110001101000000000000010000;
    mem[114] = 162'b000000000000001011111111111111100111000000000001010110111111111101100101000000000000010001000000000001000111111111111110110111000000000001000000111111111111111000;
    mem[115] = 162'b111111111011001101111111111111101001111111111111000001111111111111101000111111111110110001000000000001101010111111111101001111000000000010000101111111111111001100;
    mem[116] = 162'b000000000011001111111111111111010100111111111111110011111111111111101011111111111110000001111111111111101000000000000011000000111111111101110111000000000010000100;
    mem[117] = 162'b111111111110100001111111111110110010111111111110011110000000000001000110000000000001011110000000000001010110000000000000011010111111111111100010000000000001110001;
    mem[118] = 162'b000000000000110111000000000001110011111111111100011010111111111010100000000000000010001111000000000001000100111111111110111000000000000000000010111111111100111000;
    mem[119] = 162'b111111111100100111000000000010101111000000000000000101111111111110001010000000000000111001111111111110111011111111111111000110111111111100101111000000000000100100;
    mem[120] = 162'b000000000010100010111111111111001111111111111110101110111111111111010110111111111101010111000000000001111101111111111111001110000000000010110101111111111110100111;
    mem[121] = 162'b000000000101001011000000000010100000000000000010011100000000000111111000000000000011001101000000000010111000000000001010101010000000000110110001000000001000011100;
    mem[122] = 162'b111111111110010010000000000000000101000000000010000101111111111101010011111111111110010010111111111110101001000000000001100011000000000000010000000000000000100011;
    mem[123] = 162'b000000000010110111111111111100001001111111111101010101000000000000111101111111111100110011111111111100110111111111111101011110111111111110111100111111111101011101;
    mem[124] = 162'b000000000010111110111111111111001001111111111110110010111111111110011101000000000010110110111111111111111000111111111110110010000000000001010011000000000001010110;
    mem[125] = 162'b000000000100000111111111111110000101000000000001111100111111111110100011000000000000001110000000000000111111111111111101100010111111111111101010000000000001001111;
    mem[126] = 162'b000000000000110000111111111101100101000000000010000011111111111100100010111111111101101100111111111111011110000000000011111011111111111111110001111111111111010111;
    mem[127] = 162'b111111111110111101111111111100111001000000000000011011111111111111001001000000000011010111111111111101111011111111111101110011111111111100011101111111111100111100;
    mem[128] = 162'b000000000000010001000000000010111010000000000100011100000000000011110010000000000000000110111111111111110001111111111111111110111111111111001100111111111111110010;
    mem[129] = 162'b111111111111111010000000000000000001111111111111111010111111111111110110111111111111110111111111111111111001000000000000111001000000000000000001000000000000000001;
    mem[130] = 162'b000000000000000010111111111111111101000000000000000011111111111111110000111111111111111100111111111111111110000000000000000011111111111111111011111111111111111100;
    mem[131] = 162'b111111111111110110111111111111101111111111111111110110000000000000000011000000000000000001111111111111111100111111111111110001111111111111110101000000000000000000;
    mem[132] = 162'b000000000001010100000000000000001000111111111111101000111111111111010101000000000001000001111111111111111000000000000000100100111111111111100101111111111111110000;
    mem[133] = 162'b111111111111110110111111111111111000111111111111111100111111111111111011000000000000000111000000000000000101111111111111101110000000000001001110111111111111100011;
    mem[134] = 162'b000000000101111110000000000101010010000000000100111111000000000000001010111111111111110001111111111111110000000000000000000011111111111111111000111111111111111010;
    mem[135] = 162'b111111111111100001000000000000010101000000000001101110000000000000010011000000000000111000000000000010111011000000000000111100111111111111111011000000000011111010;
    mem[136] = 162'b000000000000000110111111111111111010111111111111111011111111111111111010000000000000000100000000000000001001000000000000000001000000000000000011111111111111111110;
    mem[137] = 162'b111111111111111110111111111111111101111111111111111011000000000000000010111111111111111100111111111111111011111111111111111110111111111111111100000000000000001000;
    mem[138] = 162'b111111111111110110111111111111111101111111111111111010000000000000010010111111111111111000111111111111111001000000000000000100111111111111110111000000000000000010;
    mem[139] = 162'b111111111111111010111111111111111101000000000000000111111111111111111011111111111111110101111111111111111011000000000000000100111111111111111100000000000000000110;
    mem[140] = 162'b000000000001011111000000000010110101000000000011101111000000000010000010111111111111101101000000000000110011111111111111110100000000000000000111111111111101110101;
    mem[141] = 162'b111111111111111011111111111111111001111111111111111100000000000000000100000000000000000000000000000000001001000000000101001111000000000010011111000000000011000011;
    mem[142] = 162'b000000000010110010000000000100110111000000000011010101111111111111111011111111111111101100111111111111110011111111111111111000111111111111111011111111111111111011;
    mem[143] = 162'b000000000001101001111111111111101110111111111111001000000000000000100100000000000000011110111111111111011001000000000001011011000000000000011101000000000010101010;
    mem[144] = 162'b111111111111111111111111111111111101000000000000000001000000000000000000000000000000000111111111111111110011111111111111111111000000000000000100000000000000000100;
    mem[145] = 162'b111111111111111101000000000000000101000000000000000011000000000000000000111111111111111011000000000000000001000000000000001010000000000000001100111111111111110111;
    mem[146] = 162'b000000000000001010000000000000000101000000000000000010000000000000001110000000000000001000000000000000000010000000000000000101111111111111111110000000000000001001;
    mem[147] = 162'b000000000000001101111111111111111000000000000000001010000000000000000000000000000000000011000000000000000000000000000000000001000000000000000001000000000000000110;
    mem[148] = 162'b111111111111111101000000000000000110111111111111110101111111111111110100111111111111110011000000000000000000111111111111111101000000000000000100000000000000000000;
    mem[149] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111101111111111111111111010111111111111110010;
    mem[150] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[151] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[152] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[153] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[154] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[155] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[156] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[157] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[158] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    mem[159] = 162'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  end
  
endmodule